// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:56 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
DK41g5fK99/nWU2/1HPekfeX1DTxGN1XwTc1anAxjBUkCfVBQh9VU1did8E77K9c
U9K4YLI7v4BfTv9fIEpNm2V6Lg4GXhqlEx2Fwp1IE6p4WwwxA5+uyx/j31AnrqzA
40pTm6ECLzrHc8hUtpnLagwYtItfiRDnFMuHtlFsuTk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 9664)
jf0Q6plUVuJMGuZhVGXxYeclmvfSjOr2Uz2NgF4ZN2Dio7vuOwgOLxQEbGyl1B26
rEpZZeboYkSPaEeuOP6fRl0r5Kj1ganN/XbqIrEsAct+WCh6PK5O8N92/gUdkXqv
00WSwShia1BeFB/5jJlPCrp3U7JA/scbLLvAGvm9lhQvrutSwdpIjOkGre2tG1Uu
YouQUGCc/TR/Z8uebIbVN6PsfTTgokLNb7NRNJWYQ8MYGv23HwBrcVKFzvROY+ns
hcTUiiAQpGlcQJOlGtueIA/RIyV0tQ+GPCEZtAIDPf5me6jn/WfFQRre6rgezLEs
8Nnk1Miwa8rEtDjKOw8c8HkSI4negacdLnLQdxkeB8PRM2kU7GUUcJKxc3dRdTiX
c2zybnTShR8byrr8+FaHnIVlVe0Ho1wgU93ZAQDc4GCeZxBtetdTT8YcHxhLcFD2
lpZHIsqcA3pV+wJHuBJSmGf3rhYJWWoIrENA0mBKCxZJkqTEN6DVu9IlKxjxnU/+
qqww6iQUEebQh0n9GF5k6WFgqvpq38FeOAhunvsEZMvnOvdEF8xwvT6Gcf+QJFVB
ppvY6HPIFsfcoLWQhGJ+XBTXfSxUoKeQeu2EZG16W0JKV31Ux5ZWJikOhUv57okj
nKcVyxJRWPSZKmO4CodJpxz6GHXA0siK5fjJ1EA+SVU8YXbqWwv+tkm4ih4/dvBZ
4V5Rl7tcnDOTyOAEnnyM97GEJoe1d5TRYU0BQNIzrgT/yFNs+SiigItPlZiX55Fj
+jghunJ7MuH8ksWje8BnCg8mvv1wdw5Z9iT6Vs3jL+ozP9pIc51tD6W2df7b0Yxj
iuisX7D8LIL2VCsJR/xI73+qMI3MmbZ0r1mC1fYKaCXBQnVUIYb/8D/VgzaoEjyQ
J+NGICriceWZ1KPii24eA8EzLDcY+DLHhJrRyk8bgrdEww7kp3gzcDvjenUj19Hi
WhP+zEv7G6BoEFXpQLPUnXPn4M6X//lIJ0eYgBJ+fEh5OyTeGf3Vbg9wXGJzLgGA
zHWa3ZGECCQtIXuHfbDfwwil/BBzGu0vD0o896R8Qh/CNNXs8bF/iRHYiR8yMGv6
gpMxMfoUT189cH9tjJWQuqrZ86HN7Fmt2xCjlmkgbhBfO/vhUbv45V9Jnsgi2RMk
2Oo8K/Zt6qi3FpvKsoWcO7QdN3WDb/E5Iaq+zgVbt4yViQgN0verN9imIMXh8pqp
aknh7B+NUCoPyiXJ9ZsJmryIAysA3i3Yl4o+MeZ9Fa5wy0RyAquv31naDBRxlHZI
Ej+ksnYokIsR7CJ5DJLyBrS5OL37IftKPSc1GAtbRHvrDnFPEmRctNPfKmaA0IKQ
MNdb5mE5gpNvUAYdBSE0QX5CzpM+OkjfwLhKHJ3J1wYDpKObHRyDtCss6/g//ota
QFhraTVkLKtmkjFX+Lmwdr7EBag6H5MnNlb7hVLNnE6BSAhaECGTIZD7iUJe8QPz
x306mftN8f6QaVy//oGydCJ8YF+6BPraey99cHudi1gUG+MXGi7rfSU7dlqKXyT/
hmleKt9iiFsiLQC2g1x0d9mKVpSL6gW0ZmK6xnttAkXVq3eRV4zAYu2HG4vV6pF3
KHPkthbAIETPT72ZTAexyoC3MI9EY04dpZi5fkcC2I/LzgGsDObydfx+FbhzKUFi
LVTRSTFoB+SUR1YfECj93Q2leMIbhdaa4bAawTEXm/rzOl4Ndk7sH5KdzR9+ufJM
jXKiytkv3aX7qj3K4evhCp+n7sjyJ/FbGdfh1Ci7OjQWik2cnH9GbrMWVa+Iyp3+
TDjdFesKPVfx9dcif+fe1hBwJ5QpC5JNY7Y3eN63TquVuzWKNg2inee2UMuMslrn
Nv8Y4Vcr5r8oog074CYE9f5Y/pkXHntSlkF8ovnF1EiiFpJ1uyJ1mRS0cjfBAZ+r
yWpII716QWkhhE+aMnn2o5fgmT6wfxWaEpPOmPkWvipC85aRahE6e0cODr/rYiHt
sQkTNRi30/1uXtFpIr4NOtFGEp/2R7/jgJ72qPFtoOjEs5fVevQnZYOdurA+Ez4S
k6nF5oFO8KzacdR60gH1HUKVpQ+4yR72hl/aPo+J+1VA32W//ez7BVo2xCiBF7yC
yDO2ZwVky49wuntwT2j462Mx34YeIfILjRlS/a8omRIBjCZrHkE9oUJ48EOR9zIc
84DrYOsbvXLuq5s/2PrAvxpAvGeo2YIVt22Yue1PnJlt9gv3fQtqFqaPLmZTEYIz
yXDSwwYifWXZDBeVx/7TsrO1OZsjFFb8r+SDLMqH1fo9S8SLRuU+QHsKVYYjOdBN
evn7HH6eNtf4ImjbiHdB6VSerg0bNGdhd4trhfO9Lw0OqBekrtG55KC62ECth/HK
pKRfVSqn5hqMkz94NbxB/yGaZ3cSd3uhHgI4c6I2Jx7OxEli4KB9sDgwhUhR1r3a
P1hWYhpuv5CD9h3U5BKtq0ds+5lY5j9B5qtr3I5/fTMZgdZJ0wg5bZBrLyf6/CNI
jQUV7fS5/rOc8Dm3yW4xJf+Ret2sXXmPiuHv9raCAtXl6KtDkfj8AJbjsLov7XKZ
uURIuQdb/g6t0XM1B+0y+KspxspKHp0uz7dbRtBsJb2uA7GS9t8teQ2XuJsiBMNx
nacfcMRcoMNZVbNJ6egKsCyt9T04fbUe++4XmQoN6cwYHqmC+U4aqXsIpNpPdrtS
XV3DVokN2SGdTjraICOe3MD4EQy/sUhCCXTLuTvLA7ll9hLhcTcmolbTZU9Ws2hi
hOXvDAFXRUiCjYO3YttFsjb6d1rq+RbXevkXcRYnQTrjceEKqN4lSpxJMwI6uLdO
CnBxft8aVD/vzjH9ig3k8crTHjpDBwIZ1yRp8n9vq0/u87Sv2Ii8ss3dCTuQspQn
cx+Qv+qpdzeysnMazFjXJliQt/LS4akQ3OLSB8sjMyJanpxXhi9qikul7pHSP+Js
nSc9BIAoCEmz0bYxTpAZTTe/iwhrseEmgDiwU5w0Zz2mU3235uVq1GUZ4r8iU5Dl
Rk+oyQniraPGEZwTJv6AcfgBCv7uQVPISFWyB4dUW9ZVA5yZuObyqiPtSapEyhsp
f43+/GrdYiDt+nS8Gh479kvlZvHrD82a8wx0zOMegDPsbLm3TYsFaNmh6RveTARG
++a7NgQ8gkEYTupPtfNbpxYS6377k1hM+bZf3tGMLNMCsvbNAtXBSfjwrmo4HFq7
9pwMWBWP+228/3MJAyulPvEIsuvjvEx2mlAPOpHNkK2yUkG61DXz9PN7k4l8ZXda
75SaOUJgDLrrcPbtqXv4HAZ4uYWfi32N9eomNAMrmDLtDZPZooNN/DBlIxgrxWy1
qAyOTkyS6pnD5TIjhDnxa66/rnhvnn188ItK68WYb5i339cAFKx5DGAYCEiQdXRY
kjYs6ykMblhAO5LcL6191zV0pSMeXbsb3XxiKtsZFyzlhezT3wSnKvhXmypIzIaY
0bDpXp7CCMv67j7LryClagxpOFcwn2BddybvNrw3RxprbdK10gZoyMLdMMDfstOO
2JBTlg4FeBYCzdoRfzbSNvr2IfiOPc+fINzzQch98bPjt/vpOYjobRG3T+vdJPnO
w1iNeGEIxBHb34YmEhtHr34/q0UYWQBXvx53llBETnDDC4mMZd0uSQPaH430UakU
wcGoPIOF1GwAP6JN4Vg2dpQk8GcTtN1MnLZn5hviBC4eU6yRR/NxnbctBrhcH3p0
iF5IOPXlwnitG41toIxau1kzxvs+9d2Jm4mYZeqxcbkGNwxIc8e/6Xllf42T7pxU
vwU0QtxX2pkwm+ONIigaoBYHZZNn5jnRSg+SRLIyltEVFh6TEfoSwP5g9kMTMSai
HRx27l3ZZxRdYY0DpjI6sb7qrwcOg4s8AzL2EMRFsHnJEeeBLkeKvTPGGsZEc70c
fyDyuUdiRLkDMifBjofQDoULw1A+CEjXkTMEPJTuA+mNKKq/eoJLwnIKuJVUiC+j
kqc1Mt0ZKPuJFY5HUaezQP/4Jj06A10Q2ShUYVxCeuqAfSHdoJh9lRMr2EntqJzh
C/Glx+noW9IDcjZAL9hjA/uX9O4MYrnznDKkt8MqemKoN+l2jdwLyN4WAp5MO+2n
pNu95KhcA5YhNVTM00U6AQ/0AnX/IafBJss17X+z6d2DiP4hP9IO6XRKlsCo838P
9ZzThDI7FAnHleUWJs2iFs2KXLqFm2OMSTl1YO89sPR7KqeHN9shtG/DalW2MqjH
HO7dtKrtbSaoRs4rSlJ+3+vkpJ3qvdUxsSiPA8o+nZoQz72cWMt5eJYIJUi//33U
7aV51WVsDsBKkwsuwWiqZAEEt+W96ZiJUSdT48A5CW/td/KA/T/pmuXG/w2Tf1P8
+rsr/0aUWzGexTEegDQthrWc+mjfBXOvXnI3Fb5PXxRLrpKwcdBHmV2G4RI6iR6D
SE2X4v7u8xPSvWNFmlojny+93LBcKZ35nPegoNxJ2U5R2JqveTtvVyIg1jEEDCpc
4/Hi4IcsH1xKpI/HV/EN0YQUma6i8TwNtiDXat97Zu1db/J7AjoOM6ggTe45F/Z2
j2uALS0qUJgJnH61AgkIfIsN1t0XiWRdJ8rsGHKWOkD0KgQqL21o1Ke0crOIKYAR
lN3Xh7RFtVGAawqGdX6WN+KsMS7zrJouHH8lJnKXsLHS59gT4/9lXXuwzqHcGvY5
rkMk/MtrWiMQ19Sg+aor/5jMOnr5hxnfKk57/3FGaWUFuETLPGk1wmRen4OfMAQl
JwiUZSN8LBO9LgYkCmjdrCtBrYQhDeKXxBH4s3J/9tnYbRwvzNHxwY8KetDpY+o1
twNlAFxQKNy6HFSxWLxkh0DoHocudpDlg/kmV14sR+EBGqZc94TuDX4wzuhPqesZ
ahfb4dO6GmlH03cor4UampeOvhaFDFvCtCPsEqvB6wGlByDNQt2h9prZ82be/DIv
qLiooM2Flccxn35vkGGFm+pszGmbiVYCPTY/E4jfTVB045NsBVSIqhkEvP7EMm8q
yVgX9GnQhRC1JrcUS192d2DCI5Z+EMejAFGIzm8rPQqBorIkEZ5jn3Fu+gh4rDQP
yTcSvK35MxqWtjNH6A4s2cBTY6IRK2TI+7SZkkSgv8OKuaBtdQgn/1jZAN/SB5at
7anRk8C/lp6Pi0L9JAskV6JYIxLwiYjopV3f4Ti60fguUJ0FVnIHu3kuBUN0zYpM
LdHD2cHeSTP/AglNa52qAZClRuow9NaCnB0TgVBCS8Ud9huaqrUT/DtrewpYyo+Y
bYHFXmYo2K9+EfSJ6Tiwiub4VVRNs6qC/2CELWjyIdtFF9mX90ItVqF+cDPgAoy1
uFpePtSdrn94Ttmcge4QcaDAOLT4DhNbqSSemCmMlL1M8znbODGQgRRVWtbHZz85
xb5FJFN0hhIT4CR/Z22SUvV+mTIg2q0WXHR0ptSEmlBJ88+O2KdgJIZx4WJyaexg
srMc+uB6YTA4tL9R33TYKaRv+0umzgC11Iw1hH9q3kg8NZU+jm12bmzfJwu5cxT3
8sSjdXSk/cYq0KZgjB6/SoWI6x/xS/BXKawomUp1CtOenMhSQAabbebf0EeI7gqJ
+SMHly7hnl19AFA7j5nN0uYCgze3owxyodUdc/9suKYIcrYJ8NJ9DvJEDOVfcs6P
z/2xGcO3X8cTPpdtruA9hsyfNWdi8q72/qfCgRIG2vEkRsmjSyQQTzNQf8IGxumj
jT+2NQhYXq1uSv6qKXY+21hZFGEF5z9U7w8oaYI3Gp9fyHxf9cQYeILlO1UaEl6W
AQxiuQlXZSigMpShv1wrn82BuJ6I2Q9XKiVoAiejsz8MBk0IZkl3LTXJB/Iytla4
FV29nUDKCM2qKI7HbBacCudUNt78aDrD+TI4vrhRHupzEzjJ1jO2Z2Ij87Du5jUx
liAn8mrweGHKxGKCKBSLeaxvXHR3UbFSvaScgYGBsaOZw/rIqDUFGiDo7E2Ef6Ac
B7ew74FurB9xR3pmewTZ3xhjPddlyoZQs0yqR2Lxl0pIIWekQc0onF87Cll+GY2B
On0SaKp68vH4HLPSRaZ3yHAmATlmCr7LlQMjw/pCu/rrojgrTpW5MKGOdk3DSjZZ
ZLkq9AU2nnjBuVW6HPasVTrm+9FTXG++H7zdDlzXtcoEpn69v4JT1HwtPiefArYJ
GItgenjZvFJg2ebp2hBG4fezVtBeap1SXgae1LLXBoimxGjA7Sz1DjAUE5YOR0uH
HVW5KP7rlT4OBernkmXnXF68phgyU2ISgpN4CruwPodnyXPGqdVFLjQYzW7GFpEo
uHlstiM8hw14vFA7Crq6pdygAIrd8N4LPsuMUhwA5yuNDfAMVdJ8tUH8AbNQkizk
kn6xJ2UNQST/9au4TrdCZYF6jqeZr+jQD5UmIPziCOyOk41l5f2MVHSL3/U+S6Ie
L6uJihMcrx1LTa4O8lCVM4paLy9XGlkbFrb2NN02hMaAVN92ps+Mh6Qhjx4ComXn
McGFzhFAm3Jz7cfrbfAjA3d2CFvJa/meWbIQOQWIHIg41UeRnpVRtbzu4KARydez
b12VCVR9nMTOw6ZjRc5pjE1OHTSmuLYEaJKoKHEYAAg1MUH4YwiSgsZb48D2quXr
AAB6Zygdtdf4vHnNv6A29bBrmeGLRb8zxtCULjgErUZiVDzftVI5Jg+BIEDqUg8B
lvJnsb9j5zEYQHcW699KLJNIior4TSCfmikarShjReJfU6Up36D7Gi+lVsQec3Ob
SD6jnx5Zr/VjXI8yXzZe+1BS/TR+jqkJZoLnZKJ9+zYv3ZwYgn0tOpS8c4TDh28X
JvPqXwpd2kzxa3gHTmi5nk47HapLdekHhPz4e26bagZ7NVl9cDJeiBa6f6MJAk//
ln8taE6D+FUjMryZsMf60yHj6GOaj27mk/vuOlzJ6gpKjT+xVHFg1T8vdmRrvN4K
X+i9SWVPGJOvH7Hf4YRKx5fhEkz7fdd4Jr3dcC25nzHFeH+PxsUlPXkyJPIeqDbs
IdpYu0GpD02vCFjhNwPqPd5IxVDuWUhfSlN1FwNcr95nKbt37hlGTvuRgtnmdxqC
VZ9hqOnF1W3ADcXaOA6Ha4+OcXcS+RotmbLvudPMEDY6hCQxu7K7jh6eIJZNB/Iu
cNlhNgmfcewGQYgDm8bEHp66F1pn3xW9QPGlgNgG9XAde1CN9BZu4CeKi9NDuoP6
OYaafXAM3MlZbRmk88LeF30g9DCh5zr4xunfWmtRO3E8F2oIZbOeAXdFCThhK4cG
byA7PrwiTwOMBmGPnJzxMXtDCOGlao7e2OPHp+Bzrpec9RTddmMJzF6Up+LOxDKf
h9QGafA97mqQrXO7dJac7FanC61WeDZe1EVDmmFwNWtoHJyrs/prKhinMX6w1Vxa
jzCmvC8clU8WIhGwnTz/pIt4S2yzFl9JWwOrok5YplU/ixdnOzcg+ubeAJfLNZWE
khtcahzBI0gqrhzza9MJRY2/I18SXdestyjCGkZHqSlOzJqcqg6V18J/PbtIjhBh
64gIsYAYSyFkCuvm8eHAulYqO9xbq23l3mHSpqOKfnE2SpJx5pC3LL18SpoioLWZ
bllyTP86Z3fBrf+OQsQII3J8khgCmWOOo+jwh1KJCqDT5VF5zsCmPzZ7vwiVNTRM
cyatyj4V/8SwjOr/oTmB7K7hM/AUyZdkQzilE+7n5KD6VAjnTBX6aSUO8OfkIo3u
uU+NcRqoiWvkMpRIEs9mvoabVf20WH+o6MwZUxKnxQ8wC03lBGOZrsBGX112ntyI
tU9iiG1igSssQWFa5LnhkhzYXK3pqmWj+PsfmnZbjaK28V3ZVcRuDQE1mCYZ8efw
6mCqXDfoCOVYj+tiNY+y3WFhLA74BlfvixG+RtQOyCA+avmkXSFtBbObsV7/Nf/p
o7LA5KG85BhcGfHsNkyO+v3SfcCpA/oaHY4oUvZJzEvDE1u2UhHSyVYsSh7O/2/2
Gy2FrjXwyXvSgnACLCizh7Gyb4/p+BsTIsWnm3uiQ0pfkygu9A+C3Oc90YT00CSh
zV5HhToMKGEILZ0LMuCv8SQacZYpVLtriUNYR4RO5rkh/LsgodtFGh/BZp4fk6fH
jvtm3wRJ7SXHnIaM8VywtavQw442xjYUY551l03dlJVcooKKPBkCroUkN4zzOOTU
Vth8gOxCLOl5FkMNgJZbB5p8vcChuj/mxukfE+0hOtUufA+gxvZgopWfRyYwOKjv
HGwj6g9j/Q/U7oq63oNTL+UiwFFTqigl1vsEZq1cfhB10atJOrA9b0Na78BBak4M
QoNfpseyxUVkHBziRhBgbh8ZQDN2DHOahuLlbTusk9uQxyFuYhi7646ybxFJPWD6
WcVivRfDNqtZM6YJcrhQvObj1URxcH/yOB0rIdbEYXFCwHm9TGPGlNEI+TbpGDUY
alKitEVRanQpdu4+pIRZV2+fGcyJ1HQaPwXANSZYWx3frCSS7ZlNecFZGUe69Psf
ZvM1THOupiJsghYtXZQ/hZEX+mx0AGY69F1r52bPh2h4NHLMTJCASbr2BpF8oGTN
Y6WNWS81NeRUYs3t0Fn1tenSkRLhgA1vc+jCZB52dWrjpybfJbAYzHYVbouukonU
hF3kLC15AaaLHWZMK4sREMONY4G4v/TjAwnb63HsvzwsJ+SYYvqQQSAKePxdAKO+
06d8PyNJFJZtiR5nmp2Lqt/QlLzUynPxFZdFyJb+yUn7jNpJdjb0p4v5CbHqDOQf
27hQwvJXIEm2k7CvrVeI/n7TA6PW/fhNG/VnX2KSYqFU+cvuiHi9GF53wV7oV8YG
daGIrqU4NUsvV91xI3g47KWkpi2lVzTqrScBZc84JwMGYlTcFrVSwf0EY1wdvjz9
xH7JH9ahI1TImoZhEnPTN4KlywuxXuSj2e+BqvMqWJ5yRhT9lI+pS5CBhxTYfZls
bchen/GLcaKffjML+XpVVkRAnCYGuhaUz1g0BUHYuhTUeFk5cs4/I5oYsvFVS0E6
sR29oBEUY3gv5zE0MI+s5r5W7DzdJsWQdS9U9nreEoNCLvQiibJ8tBmt+EbMm1JB
AZaxjjuodecQ46oDUJuePNb3hvB4Me4jrrs6TEb148QETthHPzx9MVgQf8N5LNkQ
9qiJtburJr2cIj8tYsFs5wzk4v/yy8f2cAU6vSzXeqGz7LaKy2cw/KmmPbheGEK6
/azVVeCJnU9F0m8cvvfv5DQOKQ8fTsgUe0ok3Gzwx52faYg5lMXlFlp8p8lY6lWw
Gg/X4AzqrsYkn3WYI5C/LKMfjnPg8fx1zblcOhjRo3gXQKN1DgwlGRvduxFMpNZz
xanNoDVsdP4O73t0Fd7Y77ajdU9zUJzKL/aIvpRrF8Q0pXRK7c1Mwezm18Ns3isw
LlmgEJgdtLS44tEXM5AaoY51+jgjUVcmctTXatlSZjRFj/qi+hQ8dSK6K+s3qVmB
fPh2C7Nej6NRNws3WBJAg4EKx/W1vK+uDP1UZBhMBic0usgcKaxzj0N63lowoZpL
DGvMFvyTa8+qAuyUazJCk/inpx83RGDnfUmjFlorvWzXB4fyhKQ3UCudHYAeOgkg
l6cr4LhE7iuCtb4nlACgTtnB3xB8XrnfpMXsU+4atGEUHqDKl/SZTRsQkTiyFUX1
BX25vqNTm5gZLt6aJhoBkMWYxiEs67yXb/s+fDXKN/BWSi90IJ7NRSlHz/PQquJl
DO08dWI2TfzxtyjatBbdbe7pdlH01eKt1FphiILCmyoXEOkuTjEK+gvKWrDyw0i/
P43FN2mknQwNeXd2EClBwcmniKGSrCn9SYdjofP3NQrDQsFqpva+p2r4jg+y07KE
mMr3C0vUxL/5QWP+FgYGLKd8YDvgS32ZkleTPxF0PuREy56/RVpaQGl5JxfmfxcI
gzxeZeTEbR5ORrM9fG2e+6efIbg67zpJwKO4e1vTEhWyVgKb/1MFzn7udG3IWpJr
GUx+n6kt6HaRIMzDKdaSvK8qh8ztMhLYu13wj/eaxkmlpLmpgQZBzT5kTgQXvh1m
Ay7dS9L/aGuBQk0YetazJDDtjK0h7UpFa76vqBT5vHD1fgBn4HEQLLiAvJ1LX/VU
boZoK1/uAiYm32lofYboR6MlOzb5eYkdeZVYO8cHIF5tvcAm0DDglX6sBd3AfZM/
0R1ckxvI/Xw4NazmXYNc39VNnSUis3noI+LgHEMIKICMm597TG3AXVX3j5cAV9Yy
l0ijnBlx2k2KVGSxbkNKGUja+oW0zIKJ7avMkX83zctXUzuR/CGbXRK6RJZ28kEj
tnxm+d39GSrCaSGTh6U0A+15ulRKZ5ZtiVaS14n7O1hQfhOLG18ylIvwDWnUIoYk
6aPqg8aeIIJCp2sE93EUco/AtOD+M/5+pWgDeiNuezZiB9qvbaPBspf/Y89hTVP1
eqOjm1Kyn/PRkL1dkdzFZLm7Sf56ZP827+SMDuHBP9t43V1iRbSg/Ay1Em/TGUrA
jPqOyDjrTUmsGreAGrXT29lTJzXq2FjiKmmgsjpQFNQaBbtCDaTcfIRCPZV/IYb9
Sh/sjIG3xfxfWVIhxgzu4GJGHwS+DXdc+4Y2cMk7AkUT+kDDm3xSZeEOuikdc7+d
py3QGBMNnkAE7OeBAMBlw3Lb/HX19Ag7BM9t8UkDB80zI/G49RRCoDEWavJRyn9m
r5hRsz1Zlrc55imILs21SLSvr9bQ2tmo4BShbN7DNGoiDiZE+/X1h5q9UoyNHQtt
MDYfpODtKUVmOIhiUF3CIqwKJP2uglhbhjPnz7fuhUFxnoi/2ZpkDQO7QcfMzM2m
U5uOTiZ3UuibLpRSrw7mWzxcH52d0WIkknliEn8SIGdeo3+aRQsg7L0Ci2wvJdtb
PZJf5Lw0OgiOtKU7otLdPpNcyuz9ke2Y4bFXJeRUaHK/bRc8PTEtDJ0kj1RQkTE5
7HsEwSiG8SjjsLUSRpWIWhxGIWNxHPqBJEmhwW9PTUMLO888TvKrOJUGmlsnqqSp
2u5s4avzHqn3CcL+DTz1BivFDjauQOMr4t9Tlcmm1gewfP5zLZPzqREA2nU9mUvZ
lXobE33X8S1CKcU/cM0OO/aS7gUlL4UG8OATmAkMO2WnH6Xr+QnzqtPSQMpqFsqK
AD8Ex/cx1h8MvZwvdxCq7F49M9V8r4TVVVMOn4Zyh184r7qaaXJ4VKVMGd9Iu58t
eHbLfMGXUDCrG6PPwgKPdcTQyhXZeJggbGjJXxKMwYC54RPHpYb/Vtc82mCNMHmc
n6api77Ohyd7fqbCw/ik9VKYV0ldtKpWQgBk/OnXY4dwD3vNFYZkAet0uzRjZlnw
45518QCqJBmyE3iazA0zF9clq32nvRbgOjk9qbz8jcz3tAYFPv/bWGlCUweikE1I
/VcRpX+jZjPpIYE8DHBUG62wxj10jh/y0w/wbSEWwEkGhpn0Ba5RXz8WPveFQ3nz
zgJaZTdlMj+AOGhhHstWr512kr17VMBF2qo3MqI1t0c7C90dv6FFyJXlDIfwKf5A
nVP01KMU9GOQvNfvqmNpgUQ1rgBHHlPqTKR9OlI/bD4NOmf4L9B2K/OWg92Z9SnT
MsX8RN1Ui2dltpKM9AS8F4p4wf8FinSWIZrZLe+hiX8uLpiVcBoka+++rWa3Ylfu
ImlUTPAG8RALEm+HpT5cPsTEdt04kq33oEt7l9DJrpm6LzIojyb6snMloM/f2Cw9
/2EfV49S4fKuCL/sxxlx0xPiS5JilCeqi59k0cKlksQWf3T8Vbq9DHfHyZ9VsMk8
bYoNQKLVObQy2zR802HHzxCdPt7FT7+c7g5YKEm2kniIx7C/WREKFrnfgkpr17mx
78rJWks9EVGTkFcfNt2Q7Ou3SR8+U0ZQAegmcUk8pKTYqR0pE/T5wVIEg0+mkMbO
6/iMNHH5Q/cIMlm+GZC/6RYqGOuJyHD/xj+X9IjM1DSn1w1v9pIbl/78CMgiZi7L
Xg5agE6x8ZazEuWkqhXmn1tw+1orBK+zK8CNvSOYwaO4BVpUjX7upEiS03/EdUbs
nLUGwO7VuZ+bD6bWzF1mgUevpTAvPBAD7m5t6Ws45EIoZEG4LtdQ5xZbMKyxOgj+
Qsf0MvmUA5n4gZ3oKXfx2hhrb2NPidurxhHSEXo8w00qcvgUgE+gm6ZVajaWTUOA
C+z65Fq+pgsj7nCptrC+Z5q6nyM5kxDHa/sV8NFUhag5OV65kaO/f3giOs1xAYqC
MRscWZdOYzpfwPKRPl1WpoNJSoNGs1tb0FFOea6vJkwaNFbl+hymsL5BUPZ1Gkub
PL3wNMxgBhaqmoAaGDClDcC+y4q2SHxNOjYYqzkg87Ro101IQxNRolrZYvQZdaa0
+uI2qgXFsLBP4/Vba1t1spBG3KSYZjntc2Nv0QLFiQKbT8ONl5b8eM2yOzH4DrCv
BXDmOHlLcxyi6YSabAR3+TuyNZwkr57aUmXcjTFvSRbHMv8c5OclA1V/zsK7Vij9
YJ7Jv72jM2+AlsbOixeLi98gzA5YdtJTuDNQ1RFeax3yHZY0IWP/xGjB9eb/7/98
RD6RiwN7WxEtN0Au10BuGVE3yEEfUtE4/vh36u7hdzohh502+idwzJtMHCvlWHCp
GUHb8k3IoLqKISShMHPYCUCeeBc+DIvPMsjAAoVHbxZDx+MWdggSPLn/hQ8uOJ5Y
nQ62k0JUzbQLjhZuiZ31h81pcUhr9c3EyylrqIRIEZJJ5spQ9y5HUlugUaWMX3sr
qzuHqqoWgBkDzY+8N6BHSlZ3k38tFGoHkjLi/VwTUZeQ9NdOGe8+lxksC5QDYzeb
Uan5anluz5itQRwafylbbvr+RPpgevZ3TdZKaj7PfpBd8TT+cl0/obnMcDax/iYr
mw+fEH7opv3ly4KnvJM7x8SpJvaWcufaxylbZcsiuVjPR9ip+mTr2XU9Jmszqsya
G3BuygJ+M266sdowOpqPBA==
`pragma protect end_protected
