// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:48 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
oCSa3xhy11v47i9cqZF08HiaVWWPpNdlXZJfGYSLmRrOFbdJq+ibdELAFSWHwYJA
NjhTrEXPtiSy1/cCtiYS4lEWtPPz8n+khQLHNE70VEnmEb3vVFM+ztA9w4nI58H1
aGrbkH3bg1NCAuC4VPLgB3aG/8TQuE8CNZp1mn3VVbQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6208)
5XVzvXgHSDWSeVTW6cZBm/w6oz+534IRwx66UdwIdD7QYcWkepwju3qptemL5Utq
f97tK2VMYQuEoWHC6osiHS0LrneFy84Yp59nu02GaZj9FHP3y/bEEUqJtFOi5ZKX
lK5n6NjuntFtyx8OzzYc3q+TEkvpC3a0bf9O8SfrGRTnYDEE/EaoLL3+vzuhwwe0
C/k5LNoBUVopXZo77bYTDdDFHSSdE9ePjS+AEW0W/P5A7VuMeV3s1Z12ttndo2yh
g3IWyl7w75azHvqOCUulEqRnvhyv4ZxAx3xQfhgnDMts5Gb+2iQ1aARQXvEI4MYT
hTknvSJgsMWbXIRnk5Zcvu/82lH/f5JtzM8RHfKYQfwHpfGrX1bJukcPxvpH1D9L
b4/QHQsui/XcBdklDD7LAcRQ7ylf7IZ7w/NIFwW2YQnU54+1qJm45CQmeh0jlruD
0Dr6Z5YONk6r465X71wrEZ80HzeUHGnBF+8rL3kqymwpnCfzAuavfcRdvuHDkej+
FVS/pDxAOZG4yqx0VMCnSiJ0MYZ5VugKpfLI2gIpgUyJSXolot9grzjAodhO/TRo
88vyuNpLyKuUzNxapzFcwfIg5ypxrvC8kbEcZxwNwddHgHeK9JB4PL0RUxFP6IhD
XjNVvVBEs93l5/Y5n8NYxEpQomlWzdano4RQBpAXKfRHRdYFPJ08hTqY36UX1v13
JmREPUmk5sOxlIOmI7jBWNBlmK8K4tFHb2vShkQHiIxeXj9IUePt+J/pKg9f8xDG
+kqUbAUq0Cn1yR+h9xS12ZlS8vGt/2E8mJ45WeEkRV66exEt2SmKhdgi4WkVGWTg
hTsHpyV9qh/m9r0pFj0W44PrryaVdreYz4u5r2XJHdTc9joayoLdOnoz2VKnIocy
8ysXWKf2Q5fB4EBPsLOGGiRkr/HpKZjxC0UrGY+qEBC7Eq0kAKoi4ULjaaU6Ia3U
dsLiRYWQOnOmjeQ8a3KFJp/pAEw9peckv12gwDI9fEW8erUCdPzNoa8xfrx53c58
f0jBcNj2HXl2y3eBi1nr1kdwgstzB6BHatR+6x0yEoQXO8lJKs4iE1uVUSbvjuhz
slbH/9+Kb2fNBIH/2wtoThV2XsuzfDSsUIHuJQKVyeYRVXe1dLNAVUsbk07HiaEp
GCGP9EHaHtzDp65D7aGxGln7ZukyD+yFTgCGXLt3+E2q0IpKI9TqbLXIB5dg0wGC
5xsabNRafBMk1QyfNAwXaQMWtmFSY3LASNIs7BgREYlGWF1iTu3CzkoxXPMO8JlS
kYoen8DVkHGD1f1Ff04bn6XYetowLCU6dwY8rWir5g6tye7KaxoYMTEqrBTc9CdF
TJ7Z47KNj9MV4TT74S7NOyUB7THEkiB8vcr5Vt9Kd6ab2nOmVrme8pbvIRUFiT5N
cCOvbcG/RWpqY5zLWoibk4+rQFTOAHhHfFLtro/kT7Uny4j1bQ/PvoMwFCoJ9BPS
38qrTBVCLrN/Iw5JV53YgEObkOD7Z54h4EyghlkgcbK+d2aLzVgFim+k45recHFE
1iY6r+TQrNysHe29K8wg86uXv/8sgkcsf32ddbU1nBHTOxRSVoDBQD5aSr5Sp/XK
kP1rpViTDJDWgXpH+bau9kBxJDggfBAndXvkXMXcqn1kRU7O4iYG6rYRegXEZSRL
VnAdiNzsrx3aLzKuhMP0mXvMn1LYzpfHNdA/QvrlwLr3V8vSWs/l6xbb2UqRpiBT
d8Sx1AP8Ijue6Lwo3CXfMyZFPI31Oi8NFwDFLuhEAm3V8JypuaZHW/V2U0xGUVu/
gHpKtzLtrCG40R69IlBPNVz+r/4SNrJJ+BU4YQwoTd91JTybjVDpR/9LZszmzRES
iisNVKcyYplfEidbWL40kK1xvGpaNH1AGlGZJVO529cRjY87EagTlygMpZPKXFP0
okzb7GQ4pywZQXAWweAkExGKpEBk7g9c240advFq3CgQZW63ttojY+xM939FL8Nc
5nPYGzk1/wjw+khC6NVKyhqUxLxyZp9A531lXuL4Q8etO31CUZ2aOOrADZTfNi1R
2474yZo/4fGdbe82uMM5rf793UH32tGA8s23e2CajyylojydLFp/PhbdMArMJ6TN
lNlMBxKLFTUXgIDeZ5d+H90SpFFrfIL44KE1Ds9jqtt6eDaiaDCMa6BTe/ra8kfC
EgXBjzum7xvsr3g3oimESo3+U6TXdMjdhUaUHxUQxSsZV08dWSeOW3FLouXn+ebk
g6PXdbQAdSUuqJpCijz4r1msD0QaxjO5244A7gcgAghM03DSTWNicER8skDGyC+C
lqMKlvaAbYWeNKOw3IciRQryPgalWIsxhlx+XXLu4Jzkco6v4RAzZLs2F1ICZ4Xi
KOOkEmod7DL6YLLskyTpvj37yIzoBjEBk+zXrWUMhg9xVafq+j5CVSqha6VksAnK
QUex+fQs6GxSmCfJBJMvyfj9YXTDyYJieg6lD8XYEWVoJyg7r6V+njWXx4/FogJg
NjY7uiZpligNmeBA95vHrrioMJ8ndyMAcD73UBN/RddBkieFzhM6bwoKC4JwrEGh
DjzP228nYiWqIRfoznpzajPIA8CK+r60Y7X2joZ3iFPGn4zF12EDHt9LzQquNaCM
m9XghY5ZXbiXduxP0ReYmeckqGM5SNE5b/z2rqgvITyv8oOhp6401So0xEHPGkAc
uWJP+FyuD8zdMdQK0NwcJ/VtgbB/Lhwc7Fayde7Htm4Yx08ENsUk+cLcPy89mPS+
Ti+KYvkVINIeKqUDhOGCrkEGU8fgyOB4k9Djc/b5Ax9B/o+RPV3T11ri2UhRYmxW
8uqQ4/waJJ9WCb6Dj+NQuZ/Q6Nh0ztJD46gmIbOEkMDRjCkm9huzL9pAWJ8kVv0u
DYHiwIE7JbtbK/aqom4YCQjh1LbtdlA2i3uiTGTFPcG8brdh7ZOIY/qBFJBenEdV
lQfY+KYa5kftI0gBNc/GP0g6tR5W8WQVCDvpqaEN+Tm5cN/PZ+/tKumb30RsFAwb
ajUnbnio4QUXKdqQeiZj3pdRaPzt0w1vGalhkFSVn2n3/v3vy223Mr7rHQ9eQjzf
uD0LdZ3Yl+5t5mUmcW1f+P2JAn8kQWLiu9//olIY1MiyB/1lmtrFr+ZWFbXkLb7n
MQgc1iFsFy8qqlgeKex/saVzhhVFcBkbUWIfYldk3seyL+jyaI+dQ0pfZhoYF/eH
eVEvU1x0tJU7M4HwyBg0PXjLEj5b94FOhA7jSmMiwj/et+G3+X2NErJko6k8a/Pt
++cFcp3tZiBnzNk+Y67IeaaDCPt8Fcvh43eC0iVTHJhaqYf2rsMLg3BDgHxojriz
0F4lkch9DNFbAftaxljZ7lxfrWnJjn349+5V/hC4ICDrBPBiYIdcJjERt5WgeAVV
r7OwwKZhJyk6k4NkhO+dEXKZnplRs6xqbdxPKaFhe/Q5XOKxVfHoWDTQWgDtmiCq
xCZ2tKoCC7IN8kOzpbpvGfY7rsiw+MkQzJqNt2wEHkUzU/6gv6OOvmmbeRK0wuap
gFU6GOdnPIAvo3MLUsy4h1i+rt055SptCNaz/jq4Ve4jV4hNeZA4XSLQgniyZI+v
si1jkT0D6q/N30kM2ajSpYES5CgOnmrcCy3FoL3AFbHCX6cVrATUOaw9tBewPnWt
Dsh0v9s6y1D/RM3MkDAVLh3vuaYv906PZhtVemu3nDo5RWQ8ZS4jLcMWwp7DdVof
NYYQ7c+UFKfRFYCx4hQNfS7imVx6y9Lwjn2D+cmEvu6+06iHp0/ziNTBoLgeYf48
kn4otjB+xUeu+It8hOLf4mIcguAWixi4dhWDQSKMe0fHH+2VVn4XtsneGPUI6dp4
wm1FzPKg7lM+9z/pfQgbX+wOXLdvHYKFbmueR8LwuARdfzlYTvGYm8AAycQUXw5G
xVsd//cjxAcKEM+gI9RLLQciBco+Jm2kYzUIYgqvuKu248OnUln7Vh8ebNxESbed
+lcxd4nqdwl014Qv4eD04A9fe93sWgNflpVk2L5UfnYVkKqdVxXTYx0APDOSwFDE
GNcWa+qKlxUglqURwo9W+l22pxlJPmeYt3h6XCflA2Ye3Nh5saAoJEU+YmZI4lZ2
Gyp4vq/LpUp6Bv8QKJuKP7NnrHA4eVkJ8NyyqsiWD/gF+mR45MHPmfsKuKs0WP82
IeG+XkGkPfhIfjK7VCuKeuSLSEN4CAR7jZpUaMgKRMKrXZ5An6nw/K+ZkxBBBGr4
j5EtZ9v0jMigs3anjLsJolFUgIDanE/7NGh5Br2Anmv97orR/ppeudJBt20uDydS
r8q5/jwhf1j/ZhVxzsmJU5AkHA2yioCdUCKVJJNr3++IEb4nvfSMId7YfKRhLspX
+jwCgqG1+MCWKRU69YOdZn0PlSYu64E+Ea6mH5UdXJqauxdJHwJqbEy0uEfw7MP1
+RX+iRiHLWhNybdOYJU3C1AFslvbozjctP0WLMPZg4Pr9I2GGkw0W/xwdeV065Su
L2Uf/6Yic3Bn+4pis61kNjfapERIx4xbm4YdUiN4Ycnvu5gdIdnRFV/955qYsE5h
fgpGrHqA5vj/xUg8rINLt45En1RJazvEXFMRAvUHAGIx4QY6qM+aaLqsOrdhStW+
5fTaNLTczB7N4Dg5AYntJEvVqbaK9zMurzx52MC+u2oLkrianYD7oChCdL2xU1Oy
UUCD/TIeHdNq38YcHVLJ1OWtYebQRB7t3AVUGXD0ve6oqp4L/2Ug/Q9MHUy8srDY
YvaGfoo3HM+jD7QUr4XVq+HYd0zDgNEBN+JAegxkUH3fefRlp6GGapiklYT39BDd
T0KpsFkfaI2loB1TeFyS3UR1SRsWIgetNh6eLD0vc/CVDHcyZiVc6L+BmWNhoFhp
S7Fl7A0lNRdrADDLC2oQeUJ/sVmTRVuv9pXtJzW6HDwZIQ/ls7/gUpJsX6uNaTux
FspbhTChUWARz75MfAzQS9v/4+QSTmw7Zxkzozfdd7+uvwvk+VoPGZahzp9ErNi1
sOXXpegN9xpps6uLvV1kvvbUYaGGtAifJDZFINpMf7ZXtOo1yVAwfmG8ij5XJc0I
rSTUJxClx8VoSHGyd4T8S1Vk0MKSx3JBdfOm2HVqpuDJyIL85KwbkRhtwGtpo3oO
gcCmb4ObIu0cK7IUoRNj4t3LfBrOmo5NKWPhb2QykQPcjuEBCEARRCi500YVIJFh
OaGz+GiNkI3XtfSpmOpwfX177gyahV/0cfzQqoIp2DjRHltYDcG9TwrFIADUKGI7
iXNssZEpkh5KpVGBMZlL/TNJDQoY3vj0plJjdRx738/NSyvMorFo8omK38XJv1Dz
0TE0tUv5s0NFwj+W3PkUWw7miqbSvdOPBwHPPz0tsXoAR0or8OcyP84Jc/VRM3Yf
EVWrx1pV9+cqCoaWVUCISIhIBtCdNrsMxfACdPaBDgTgcv7hEqeyUK5BN2YSjQdj
nY61SuKDa91ErOlufyopKm74sKTlZbC3EZsRPYfGSvU0wO+doe7PniMGsN7/3qA7
WFXxhew+SKcDXJJ87CXSmZ9VKki2VNmpe8T/LMY5nO6EOW1gLA89RaubyiyeGdyB
QhPXLpYVtPfHfbH5V3Z/MERxhifTkJBGbx7DAqTApULaWAh8Q0orTMn83XW7CfU3
fqap4WoennxvxFmBWryrabehk+ds1exqVOqVloHtUsR5X5Dxjpb1FC0nngrU/j6p
OGEVgxgG5u1K0dphIQ6BWIlXI5L1k6GN3/SRFv89u8gq+japxl5PRFMG8T6LxsJ4
ysEQ9WQTyIDQzLn9f05Mk/CuPwmKuvEUoin7ACmVRhZSrR+UM04oEPE2uAmh8Qpx
fuc2XilTySyNjlht6y4BO6bPM6YGfLfmhGx+4hQVV5b77MOWLIqlNzwrzM9XJvBv
DyGUPvYd4iToCCHt680l2CoOS24Hsg6SWcmSwBIfarzs435n1Jh6q6Jhrze0T/yE
r2h0M0GqyaAk2M3vIessfZcvcIedyvGbU8a6FO7Xzl7pcs2GW7y8XKKK3UEJRmKo
67QA0yg5QEd7x60eC3QCRHlQ9da/M8CWvYLOKQfNo+Og2u9owmo5E3Xr3a/KoybM
2WV9D3vDMuabpD5kCmEMSIp03h5qargjoA+ELlSDygollpmxDvulcx0NRhLR7qGQ
Xey+ifbfBP6sOdjbzbikP13961CE3s0chfIQ7y187a1Wy4T/V/fFaY0YgqBxUImM
JdofZVKfG25hHS8JXAjLKe3Tk+cTuKx5hW+tGUYM+VS8z+MeZm40wsA4Ugr21uEM
uBpIaXCJXUYGPvyrjzQPu9iP+R+rAWVjKoSGkTtx3VDYp/oqPRgshK3M2BpA3f5Z
LAZo3jNhyVT1ceKHNnt7E3+I0ZZsBL5E3YmKo3IamIeaaG/NIQ+TPdN7FO363U0H
6nGum0CvLn4pBqOr60KhBOeBTtBso7VCYIWsX+++uG1gr33gsQuFaqay0HQ1n38q
hBAonvkCmqWdnlKsFwBfec/8RmbgzfL0zHkfrQ8nLw8BTgB8rfdXPOSQImn8px3e
IJ+ecL+jemimLGIgAm9odicpG27H7GD9du9srke6FiI1MZ3lWh1nwx2YueVUzgA5
rXP5rQfF2nux6kKNmEFE8tD8+zO5mfJdSho3yBsqyRu7Qktw3D/fIEJxrBzeUlIe
1xLWeVlhxDzOA7gwGYupSXGgytIwtmMPFYilKvgtZp7rzPgvdfrZBHCAV0nNX2He
0T5oE6qEYX8xF8Iu3X0mWxP2+MkpxQHeROW3s4d4zLQf0gc89WmCAWQRYvnm7r+E
QXrH8kQj4BjCupKMsviBNJu67Iw0yUKPNzEtHGopv4eW+3ad5O4xfQNIjWZeLSC7
HCaH+JFR3CXNaCpZ4AHKTWVCDwNUgl2Wuq+vGEZGGE+LkInQngoV62ECwMPsmK2+
HMA+zPYR+GMvU+jcMSd7trtxMxBn2fE37XhQE4gK2kL4TfdkYw0NxxxjhxleXRpw
1IfhM4Da6gu3peCAthda3grULHJurmTgCUQo+y6SSGPflVWgw+/IellLmZLbLNuF
X6qT5SRgeB+YIVRoqV421ZG/iFfxGMjrWbwDA8wWXQ9XW6/jGxORtuoZvsIY8mS8
S9/NlOFH8FCNVNolfjgDvlgusw5YN3fY5uPhqj5T8iYyNJjRLXxtZAY/87EY1ePB
ARN/F3HaEdaw7t9ZBTENcfXsDX8BKeQKiI6LIXcvvdtN7MYiBLpjXvw9KmOMlgFp
JCDW1n9Xhfj2/UkEJfBlsyLHbxTfWFXLqMbSoJ4/5xaAmd5kxGukAntF3NlV/229
Q+XNmNaXXiTrhyNGirQlg55qtIkimIMQtg5vHF9Y+sT6XTUBmaRepvJVdyl4+zkR
5SQwyvYPiTfMHJcf6PLhKg/ger73dzB71le2kP0uFwi2+0LZhSTfy9u/MwGWSQEW
ixxvRy/vuUns+VElKoUshDYiNGSfpdxGj0+BQhKFaL3mhRyNc/momAzFt+mklmts
9KBJo61/whZHVFoG1LGEep4hh/spCo6V0AJQXQB8kxxkYKCa4MEq88RGaa10clzE
FoSj/PLBoPBiMh5MFr2+L54UP2aT4iVSn1wHq8hY/zFEuixFCFgq/p0TIRtdo8of
3A9tjbMtjnkhmjQh3ULjcrWrUhyQyYE04C6yuRWiLZzhDtXp9oXCF7/zmHHJTPnI
A13gDRFfCp+GB1yLdFQxuk8ubiIf1VKCbD1vONsNgKfDeOYaKh10w4AKzn7NmF2k
6LaoAkd4jWgQHeg8n4blNMH9iOMeKhKUrw1AXkGDUewjnm8JnF/aVlwPmPyiCBc6
B9Ip2VTA9/cLcm9DU3uCQtEMSx8EGGGwuMuZBoVnXjOXHPeICQ3w7npUBXMyhdHt
QvrBhO9XEmt+as4AYfM70/RG+OFSWxsa1NmmxDTHmRcjLM+HE6lSPylREdldTeAt
QAroT0UwSNt9vR06tH4vPjapucu2FERt5I71a7zFEYp+2SmXcBQKRggf1bsG3lAq
bniLTXSjZf6HAQMS0/rJsD/GuwV/FvYDCBUj4DIkEkjwtmCPwcXrKTbatle3oJ5B
ycNfGZNXm5NtAxlS01SV4wQX/qE0mfS4lS0W6vIuHVz9rWdmv3CXCbJ3ykkmGmlW
8YoahiYPMBpkS0q5fTYdqsxV2LKG7HDjE5fRnwjSffGIh3QkC0EQyDOYAt+IS4E9
2aNqfSwzScr6wXbzPmIu4y3qzK2WG2D2HmCkfEoHZO03+m2AybPjG/eY7rU5CI/X
k2B2D27Q7gjr3LYwKuGjhA==
`pragma protect end_protected
