// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:59 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
kv3l0FjnNZ8mZHq3l8jeV63zGwKVgqWJbPmEvKtG9hilH/4cwpQbY+ZKYvf+8Jtg
6mNJ2qftSX/nI566T9sWj9TXkweKVzUhFXh9PWRFhpFTXctkkFDwsHA5YtVIOGFq
U64zTMjpldB4p5HOcSKw/ZJ+Pnh0BWpwzPZXZxc93UA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3120)
SoHJVFE+cjGXNs+rPM/z1pi1Kf8Ylpl8tvgRgmpPqngwqfusNSMGcEcfQsQy1Gfi
SO9bt9KObpwF5qicKFdL+0wcDTttTXoT4y6MfdOEZ4rWHywcUBrJdNvZlRsP3JCc
nLAaQqRfg3SD4nJfNIj5yEVK1tRepDhlCdJ9R/d6T1EE4wR3XHlD0F+abUaT5ZA4
GbhD89jpsR9fDzEI9lb7t/l8wstHkpiDFLqo+9sda9kkqnWE6NwFGXV1D/+X+BMf
LciVhpIqauYB4Y4IB2ekyokFOgwyTOO0yl/sMow4M9iTfrkynIIWM+1kkWtBYGZh
BWWzaWN5hpsUJPUb6NRk3qOh05wILBuewald1jiox7dNKoZt/5LYf16av/ao//A1
sigJubjCZ9EKvZEkzUflbS3edShuoGuvMd2J/bbWOuqca0dbL3gDP15xdGOrkMF8
JUP2rSUKlwoF+qsRq0EdPBbD5uFcHCgFbdo0rRlbAPgTtmOPyFblOh6xA4tF5Y+d
lxy3tKQB8VYKLkY9aBS0Z3T/9dTInqsJZdLjoVFi1JPiiPsHuGNiu61IJZ9ErbZ0
FP9Ew9tS6Yra2ckTXqU6dEal4Vb4PUXeV3iLoC7rhBgCjV+gRDUO2cduVDHipolx
A62f78hiAlg8CaszQv/xEuBBmXFqzUDozgjb1YKOqTQVTaxALe7S5mBdFfGyZbp/
hvwLcnjZXYwSVfaNLPDj2igt1ctM0FZeDxrN63kNHtxulxCtYdhEWQ0htfh7Nbrs
7926PhWQlIviTZiCCm8Pbphv0Xz4L80wjaZ1N8hitGCsMhZt6s8JcW6h+jf+duXn
dbLPm4jrWE6HWp//5rAVH09wo1KEnlCbhHideSQXwubSWgCdINndbydLQNA/YA8d
8LJiDP/q5QMVLmDR7x2llLUb76socMJ8k2Te69wFeF9shA9HP6KyFczlLEeBb0f/
+tgZWCpyECnefEAdju6cxWg9zScFOybII+E1p7SIMJxF44aO1aeSEfVP9EKAcia+
uD3CjZWn7gf8EOwSUfZjKc+BT8vK6DC9QraB6Sre/u3yweQckyzUcB22RUpDNKMS
uTcFQimUIcff/DT4l8RXJod/FkdhFQOCts6+Ah55c/WpmkesiF+e/L5qhaR3cuhp
KqmYd51l/inIiuxQIoyf6QO/EY5aguJOKYRXoIT/cYVtKOyEpjUMPc3Yk0M7eYQ8
YIiORNe60IR4zHQKQGldZDus/Np+xGNnqW/o5PrUfpe40u89VQQG7FJOY0QEF+GK
V/GVagKGGwNw//mkWXYX4zkuSMY0YvQ5fV3gBdJ20nSY1EqkRsLazTCBmXX18tcN
OCcTPyACPgw/X/kMeY/aEdk+qePAyQeu5xDlIFpIN9/t/oEXN+E9LB91Vuv4VJ1f
mVWZBCKasDUsYKqNoi/H4qglqEuig9ey61qU76UW3ik+87BEBgx0J4uTzN0NGLKG
RhmsnTpLD2KWp+GFgfqXzQizmOGbroJAgUzLFK5VOShmUexQ/vH6B9+VBWnyjErB
r2/XocQNuSv16t1WtOQuw80Zlg16g1KOzl+lAhg8FLUuXTHpFC9e5FhL0ik5G5J2
PF7ticxWZe/vE6hlUVBe3gUlckP+Px5u4Kkf58CA4tsR4A7C3VeY1VQUR7xlbl+m
cT+ygyP4Mnvb4TL6SoYCktcsyTmDRZqrvVOFpUjXpMDk5/aNTTZ5K37mOOE/0ze0
t4ONKNQIicZqUzX8eUQGG3DUMIFj1khemRz7a455sLYM31AdhCIbDZtwDZ7mAKIU
opMQD9mzzkZU3+IPIiFoVJ0IMXLALYbsITxAqCK9iplmX1usKe5gskGvkLwCXzR7
WYR2q/NDKk42m/wqjPDnqLQRjJHc6X1nujFvyIunF0684qNFekNgzKYfGipcIdi0
NDQx+4deHbI5BhhmkuEEP4+gokQdFufdXDXFLTHi1YbPXgtL+GGZmQ6ZuQ1cvyU7
Z3LeYs+/bFiMzYfpS71uTzq/7k/90hQZeIi/8Yj3lpNO3Iu/YE/8wF56ijMlNZUx
s9v8w8FYfrhGP5nKmOvcbagaNOKmyDNsN5l9iB07j88+yQV/q/MqXSXlk7I3vTim
qqlZd9uGLx04gWOlpTp8A5OTJiLverLa2iOS+d4OPpJ1X7QxCuPRIWR1ZpOXWugB
21ASRVJLfUPN3kDVLC7/UN3xQgOwdrN6HL4CemIKmsPAy0ilZqLGWuOPghZqw5wF
WY9jXRTw7J6PAtUUoREaM3u+/+/C2OmfCUqXJCLN66+o8nCgY4Wbbh4A0ZCtGUTf
jFSmWVYUJDx44+fId/evvldgsWYxFiadfAnDmrph68+WA7omSBzReNDtk83LuhMs
rREwzonF1uSHuCtHpnfbUtRUIQGx9tIg4qouZDSvl816ewil9GfY8j177IvEGYUV
0Tfj/ZiZIKmv+XCb7tkuaWYru596HGM+mdzSvAqv7BLuuPK20Bfx3fZY00gGqP1N
UNYKOTxchd3CGlxQd+PLXPty6sqol/GA7dj5N332XS23UdTcbwm9k9k9rxhdmrHE
qcT/1NdRaqpHbvirmknXW7zalsLygcDubRRjGMKYTeQDJb7TxSqHkZA18plHq5ad
CWXgaHV3C73D0HHgi+wGEaac0i2n5HgaHcMsg7UZ5g2SUXeynz7SF/7+eVPXa0+S
FbQBTnA7CXrc5bmZKZUlJax+yfNT61400esXpSCk8owe0m84+lJ2utBZ1eyWl/fi
KHa3TxVCyYgQFvkS0Bom0EcZSp1jLcYHAV11RNnt9GI2T7R/uZjK2ddea0kpYMbi
zX/mJIdfKV2krhNnO6NuP76gQnPz3UxJKX7+C9ojzjTzTO+dwTCgcKUSg+INVWLd
aF66j5VVqU+oq0q/eCWLty3PntBIGBRiq+0MhKm6n4u4CRRuOaLQfdojmcvYlytG
frkPV0n1Zoi0P+3SqpAvdxCOePn85kCCsj3IFI8+rhN8w4o+swOqVbfbN4NPGC3Y
G8ZF8MiENHM/nbHHnJMyZW3YVG104M/e3oZNYI+VmPRVKkefuwxhClhS0cREW6tv
UM2gmwBJkg1TJa8wCTrXwMXFwC/GWKlPcXhosJb69EIQuq0W5FRxsV/5Ks6lfoZe
y0OHCa2sbFCZKhppO58dN1HnbSUsV8gbnL83MIVgwcsdjohLP8H2vSzVm6fE7BhS
cLMHX+q8lLCyEJieRyayn6lSv7tMfIuZ067JQ4koONaQazd+VmrDJA6ykPaKVg2u
QEVWPGN8y6QIvUdh1J+yJ7sy86pNcJczZqJHW6c+F3NTDSPE/uoxlMHoi/+t/Prv
O5F0EnI4W7Yt0RM37HY1FNqcyCys1n6oUUU0Q9NSuFtGxGd1/K+Z/njPZOsS4ugL
ehNPOnUHDpAZOLtfGSs/KptYPIfrYQIU7M/CNNq2/MWMSZK37F2H5ABgsCrcUKCR
lo7bEvHE8fPUXgT1HbdGuJT7Ux5O1r3cekUyhR/TsHgF1K2evT/R8bIOItIq4jTs
YTZFn5EuMFe4qR/ox9uqShzZ+Yd8r2HtptINVkCg2vSfUR3fZlbK4tM1RuWaXchd
4dT8vx982K5uVAZW1lPx6sOCII6i6mVmOhcZTgsmvtKazWOqrNEl6s6eVROdiXob
tGtABj2eZEOC8130kf1rWVKJLcwVuumBjLiRUR19nX8lqMfpmjJ9pw253oCCquQC
WCVaPm3wiA2bfWGBabEjXmIivgp149iTfK8CA0louJvqJNsEWdGQEZVFKQIB04Ka
EXwivmTsk3CdIKJiGGugsOSGYJJ9FFuHB+RYwIdaxZCLruG+yxxT5En5AdCbnERk
gRXDmH7OWGxtH/7gUvcSVdFwqiy1bW8AGrvtXfxsnuydWjawxlmCmpcf2i+vCsF1
9t00WbMxzOsdrgpSgbMiPOAJ1tClTi4L75Pz2izpVNkjOvouWEgTkRoO24wJAP+6
BrR93qrFer6pvjmOdZ5xrZJILc6SRiH70xMio4LDmQHXy3YwN8p/qTUuFL4F0UmJ
zAlJQhixEnZGl5/OcekAj4utZQMk95ULLF2wcz2Ym+7Y03j6PCHpDtSlXhiKSTkR
AybRuLdjnSraKdX8w9bYYzNM3uYRVzSPjqLi0b1GM44xc+kNSHYbmlE6Q++31gkm
`pragma protect end_protected
