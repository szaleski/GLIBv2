// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:49 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
PS65AB7q4tz2N4DhVTYoSoZrGDXyAh4AdaG+T7GFm5C7bKoo6wxujhmf0ZAN4081
nFTSmQ96Crfqejopfa35JkIpJGEst4iHRyW8y9suXCzVGYg6tGHl0MboWRpcoIaj
9pqGQq6RTkwHnbTlluqRqgJehhIWDHMU1NMBZRdWuVY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5312)
vw4relK8WNktvqIRWceM8PGRqtZlf8fHwC6c9WTABJrC0dFWV3DvGZF4YNn9Q8O6
7pBJ4dDuLPPrfcDa/rEhamvo2ddbHkrEWIOk8rVBVVItZQk4Duz/gzYyb+9ZUAG4
iA886yeytGwBdPqZrPKFWEFWX0dbzMqgaZyUEprLA1ULtjHywHHzMoSk5wmSjDqM
QAfoL+g39rUzZcv5Mr23P+qlpMbnZ/H564Rl0gCyEDDpz2c6LMJ72zvEcFS1uE5a
J9JeY3n8z2qfAHlXDZKSDLlas4jEr5hKRyjvlnvS0fgAlzfkhxSXDP2XdBJNIrLm
9+tO0pktHc+ikzbNR+M0Cu73ig5baKcM1Nj8DxH8p93deVFxLf4tZELGneOH1Qo6
esQpKev5mEURAj3/EcfQw1GDEH7RoUxM5PH/bflqXnEfHb7GgQ4/XurxvKTC4Kpj
bfcUCyq1Xz00K/yTd9oa+EzjJXVCxVxgKbtyOJt9OAAy60E559aRJ4C412ZXI81T
hpce1TrMzVq62NqpDREPMXIcr0i9viv+lA5rjXw+nlxUolNUVmKkSi3Cb0lKJp39
1CcFftrIdcwuBhg4Bnufsvhl0l35Y66vzmUlS6RrCn23ruJjAuWNnynxK6dh3Dsa
MkGImLw5EIXJIUVdv1TsQ8tZTxtQ290ZVi60lX2aHm4WN6sU1PuAhgbD12PiS56L
lL/odh/FlZb3YhBRRpunKYGwgmDFh2PAq5Um3dWreAka0bZB+h95WdLCQdo8naZf
wrjLiTv2SC44Yu5yelkOCStIb6CEZ63U8g/zPp4Jwv/U6lwgKKmMSsWI6TBpbz9/
2w0JAuBisqX2enw61HpEvR4sN1AGh7eUv5TjJA6UD1JDvYVRQ+6gUXC9VLJAu2as
vq2d6zVyOfV9qref4ChrVc16nTUc+BBuW8j5sZx82EkFCfR78s9dHidU8z9zlEa0
Vg+dE1tmjjnJZ3x+45cWgHDgwnj2EkeTeS7aVRbl4TXVMxX2gmaZnBq1s/Cf7/3C
9I2iXu8wlT5dUKdmzH5cWiRwjtIFoWcwvePQylemO0JqgVJHdIIdZTBLdRUSklRE
jS2AxzXUdDo12Ls2YnfAr1ic2e+32/SgI8K9AwFp9QFad9J/wN+DIA05ch5kzU6H
FObmP910IoJHV+QHaoBdL7ygjVES5HZetZw2HLwbQJ4zwQaVXE51W/rTWK/oTM/w
eP9tp1Ky4wt47CbvMxsild4dEZunSWwEzOVUbplFpFQ2XnSXNKweiS1rmwnhIlSq
lGx0Pwg4FYavbP08y5RM5C72cnRVSZGhv81ph+kJQyQeG9xX/g88XGnMRGNCTELA
4o9soPEAhOd8f1uUqFgyTNQ3U47bTfoXvI3PxgFVZYAMVjb6E/Qe/cKsZ3RqWhbn
RAgcKDVbPrqNKJnuLrAgKpB1JUqx5HoaV8aQ3DfgW8TDYwQShFUobyB6EBJkc/Sc
ju05Rwk+WzsdCz/WsmphIPd6KjzGQTPmyXJc175/12NfMa40l7MZhkVZIirnfBpe
puD+jufLNodfIgB6Nv4T2G/RSV8Ys1ni7FcumlUn5RS5QFhuYzLBaAorejvG7qJM
D2TPfJVA7pm4842iUD6s7KzFNVElE5TAGBeGcAHBhuebgbJt/lSj8aZuvLkoPm2A
MQAaePs3gP8Q5Fj6/uWaQJlcJ7ai1tv550BNDQldN9iYDihMVKkiFQ1xP3Ji6e0l
mr4c+rgoSrst5/tsJVZb2WQAK0q4msaqS3cVfXG6zfmpbSV5COdjqjX1fhDkrKTI
I1qVl75LF0+IepD+XXEAEsLZMdu3iGnS0++f/B3Ox3ZNcHm3G9p0P+sdbDn51Ce0
jSdifl3wzMkQKRaf9E431PohLJd+wZTQ2gOzsUQ8/PG8PlHvhLe3DZiQL5lDdBcH
xU+OZ42lk46qmY0I7f173U83XfP0xxS7DHnIGk9rC7iIQjxEz3UGMjjO7qTC9Gcp
3nDTJ6GNh7jRhm9q7QRJrhh4oaw+6oF9HfiRSF2p8CqBrr4/OBPdIgoivtzGIvyG
n/o9b+/MfZK8hAGqBQ86SfreIp2fQ73tcWX+A9laKgsTiVhXgshhfom7KBbXKpwt
lR6Y8bqUCMuwHwxkriLvwN1LY5WEaO9Et7tbQE/K0qlK9mJH3vgNHJkWCLQjYryX
D9eCW1/jKckXZaYktaanVMHTqqrOxmrgrRRhk1eN5DXxyW9VjaE/HDXon9yJ9vH3
4PrHIMM8C87sF17D5M1eshgZBDy0GWeUrX+cH4GJ0q3meH6HcLtqaEku5QJfE6G3
qQItShN8dwzkQp2bS9fG/q+IVSELS9rzytTi64eHSfJusdU5HYnOOxRgoUQAVCXt
PP6AljaMfD682S69UFU6nH+bfBIhbk4MxKU48Ud1cnGSLqVU5N4Qm72ujFAcN9lU
Lw1as79sxIa+orkJmbTwZcU/9bM4lYBerzJdHAsbiwTOoelF7H4iZ5wn76/XR8bh
aOINQ0RAz4HUA7chYjus72eYgssL9AZ/msXgJjX5WxL5Ea+dY4gi/fd6b67DHFvB
rlKtCxd5X0BMuXqwf5eS/UQCnTO4XGucckw2GD5chZc5KZNX3EuhI4H5Y/+UFEWr
T17ox4+KdMkZSEj+yUD4JsT4huEWgksPY7bRl1+VlBBpxbDmRqrP7bCDUYXJ8omB
hv1BqQLfZ5y3gGg7WPwd3oOowHd3cW6n0EQc5dchicm23wyRwdAhkO4z5c+oq782
A6286wHoXFGulNA1YTEfuRLYlee0C3xabLm9Nh3j0CHfKmaA4Vflot4X7LhxAud9
9wbtjisFq6LTbbHMJDIu9VdRb+PDyTcSoV6GGR3aWrPa5SkwptsXMv1gpQ6N42Q0
AwNmziWcww1vyoAQbSlcta2Q915Trwvo+40n6P7/KgI4SID4EI1VzuWaxvnRxwYp
K00tCYqzP12L0FImVK0Ed9J9aj1/f50/YCt4HwlysBUb3WAQQ05mjnWG4CHhgnV9
mcY/vFGq+TN4EtRKyDIn1qObCcLi9lWAez4o0PS3mSPv+YFQF/35G85M5qThvtyP
HAtRyBSbzm6dMDhh0Js98yWIHoOR0p+IS/xJ+DLJu/+UmwCeRozxMFj2NJsSeg3z
LHlimRn5l1+OobV3/KgTkJc8PknNSyn9sfVuVdeb7VHi+sbJ51e/I46rlAi/Vdd0
7XrVGdBkanG7k7AneoZHMNnIqXeDJwbFV3jG/FEArHix6WJ27v5+BtLWGoTnvrIx
a9voDbg0wyxuklVKqk0X3+5QKCrCLVDfU0rnKprpCRCCj6oGFvwASHYe121d5rDC
dxQG36iu4s3XrCx1uvNR9NwPWvZaV+yD09o3Cdyyoj5qZxSOQtMKwwcNUZEHUazf
klFwp4lnAARMdpBuSZeOByaBGgLKVtI5tnaTAkkxAtg4HUCj42A7dUQgDK5kdcxP
6ckwsU814UDfTbX/95Eau0ukJICgtwiO3ukiZalkmvHkQUNT4cUuNtDJEuyNdep3
OMaunO2pB1tQ+UJaEMQzoPI/2461x3ci6J6DOnlJ6GmvD0ggzAMml4xDkE5pJGXZ
G3MPxhSRsGmbWTTTJDth2cM4/qHQgH9dhg8cpvA9fIQheUulMgkFEy06BI54qm2P
7ZOjHYd1y49Z722ETuWUFfQ5h0KaJxFugHWesuCEDlBntmWiBAmuTWuX9nGPBQaG
LnKsmUIyZ7ZK2rCxuUHAFBqoNyJjFVfhbgdHSSNdR3RQ5xF2wRcFkqnj8YhSWUpM
/PoBWMjcLm3M48S8CjoO2DrvUfzO/DPuc1Ccm+AdxaZ9ebGvRCRvJw3ovD2fDhBU
IRl95Y+MrukJUMjV36qbJFx2kuviBp9IDJ9/Pmwki5PTX1L9Mv14UL7pAvjZ10uv
fhfZ16FNNRXo2Q/r62OqIB4AcG0qJEak2qJkf9eoxtzcmj3Rsm9bxP1wRgu29Exx
eEooAgfnsFjnyD3AfWZ5WdzkVBG4/M+/aN+0fQo7o1A5fuu9brn1MGpl87T9kJuc
jhTodMfZTbp7U32e5IFQ9z9Mzmb0qiEJSq2Q3uA0NDxh8IUkscjkUQpv/I1T9qYo
EHej4jWdZ/tIK2cgbQH2fU5In1qQZyD3qumqvJ6X74eQSbdJjp/aqkxsOb2MywOY
ObTLjI0lyf5jqaWztNzsrheOo/LZPc6+dsnvyS5muLb5GC2WdfLRe+xOhKk2beV4
N50FM5ViaDl1+lEhH2Ux+Bj9HxN84iBKkGlk54bw4df5vbE8FS+82OJFD2omQA1v
NgqtTsKELTPAjyAXJwhWhlUffhYwBogmqFf+UhgKQ5r/1SoxGVEzByl/trOeb7cr
wb/Hw0qEjQZarvx+iRy613kKYadSxuBfDT/rRHDEZzAqops6hC9RAW6/tiU70J6X
txR7p+97QU+wu5ad3uQpxNLy5DOTQByCV+GR9ZPJ2lB0F76Y/GCXbhroGupHifpx
NV9DUEAC4XM5KIUs2i/C/Uq2BbHvNsWy671tB69rNkAp9lpv7QfIKK/76b/aqC1Y
p0iqCXln5o7eTEmOOeY5Kcyvi+rRTmrOX8SZO63vLIVszPYOao/VA5sUm8GEItXJ
0/YV/Q7TQ4gZb6EJwba1FidVHVFCZTZDrQupUyddJBHt/aqoMqi+SDx6MKkA89wl
a8LcAQNrXHZrlDISRvgKwlb8vRphE1eZZp+VVdFcOd/PqlBZtQFMw6odpTMTuvb5
BCtJRiNsVopBH8d2LchRlD8hwqNhvK/w/cjBLndG0ONTN5M0aEeEiEL8/lPc6lhu
BoZLtBEJ0925A/xrtAgh+GXX8pPpuOs76KZyUCwDWcFqjJRpkC+F/ccs/tZyIs4q
CSqokkHlo9RkZHOlJ6MnJdtmnEQezf18I6pa6GaysZHaoJ+M8efWyemtDUTi3i5W
cG56Vh14BNH2+kanWczNhv/gQ8iuWLUP9AlWnGUaCWFrz+S8wI3DMGaSzGNXYV0a
3Yby6gFxX7EsTb/wUA111hbZadvf6P8Vrfk9y6vDDnsNrJ/HGOoVxdO18Ism/v0i
yJeLGyHzxBkWU4i34/9DxIKZQM2uVnUVbTNhaZSnqeMznKM/b0DtlcXx3pDEtnr5
h1sz4Xw6eGq3kRYyg81hlxn2xCK3Lx2fo9TKs9pKMPLQhNM08l2dE0GzAyrI4ETq
usbjTQ1IX6S9L7WJpMZdaZkKizV5bYa5W8w1v9zmMIfbXg6fBuqjpvqTiIQ3oPny
NPGrqfVwlFio84UYP+pPcfy2HD/V2dPu8C+ED1Y3rYyxcSZxWphF7ep7oeflrwS/
7M73MgTPaIlO4G+b4x6KoTjZklXFjQcTFckNqhNonmGkYP4lTOMeCE6v8crwh/SX
aq/KRpKaT7rBG3HaCh6jJiKZ7Lvtj3RmrIkIB1/obIAjv/5fWhZ0LbfYLJkWKSOy
+bCqIGFPlhRhBdE2vd3XQ/ktXcEfw78Omlwz75nP0wUDEQE6x1VYqyBx5nVadbjo
8RujSZx+JrO2AkP/eRG1/GFWjxPQCwiNKLRLwLLcQdiD80fo5XxiU+1Unv0Po7ur
LZOZ4jSVNTaYHBN7nKt1xU/R+FRa/M11TuGmKkruR5zRgRhkikK+XMGr2orXbJM9
E5amuqcrw+fEPdbX9RN5kCRPlfgEVKydJIDMePI/Q9k+yIhT/kQwcd4dVpwARzfI
KyXQHkmfr0JqI36jwZXuQQHDQdsyOwQRHDj3cnhx52OKYD+iJAP4IySUrY8PCp63
gRB9DGW/FWQRAPmF9c5gaOZ2NvNE3CZs5c5+a/bxgTWxbdrKBBXRHHyfeSKYmhmQ
CjQmLyX4GgFlgAToOPzzxFPJEgrLMuFdUjJx2HyknrzbfrsQUTFgED0GRzYmB2jp
beHNzQfiu1H654FuwHHV0g9rMcWiEYbmgYe04+TnygyrFj2cexSfY/8Idr4XWRu+
46J4+jW509uS5oB/iE9bSdbaz3rT9XAgcgZtKbcGIzkOKcxIOGS0u0V+auu62SRs
wqu57vDbvE9AHbN/COFHDyx8w4x0q7qgexFaYBakWSru2zQ0HLFCpPuC0sLhfiRs
2AMdhwJ1RZYre79Zv7vXGHO3O3TBk0MsRk01Cecn10zPTidjcljfd5xIzIvblijJ
nlY64jwVIkTYlPPG+kh5ZqMHfynp0CAl5kK/of5Bx5PNvoTdytI7uI8zVJcifFBa
z0S7VPcjyBHamFtdsstDwHFk16Af1lGCAkOmRqNG75jfzwYoCkb3czfHeGTAmqhA
aQ9n3LwF5c2C7Gyv2VTPBdSrFJaS9XHBRGMlA7FBMxW9jTerhHeavpdKXqFdaU1n
KTdeC3c55jswNP/e4KJtxRU+NmkzEgIZIUPOzk0tZxXgUiPvnf8v1yXMljPBLpWh
ThUNvqNv76vjk2Zf83ous4H0iGUv1Fc1ls6mHNL/F4whSDTYF22S2mbMy6x+peli
tD/eor+hYbkS7faHhzfzgRqNcbvAkEDR2f8GOCA7psGyDVDWGu6Vh0HUN1Wo0Bpu
ymreos9CuILwA5Q7PjBB55+SA37/bgnH6MHhg4+f0inEbozKmdZxr4U23t5tA+hT
+qJn4Xnm81UCZ82DjW9bqaVKLgvMuDeaPg9NE8+3xSf6SA08vIICLMPQab8ehgF0
eRlX7eAdsz8EzABX0e89wL0EbOZJqVHDywwU3U+RZYEF1zYde/gRXMTTpSqWExbn
ctBKze2fwolOiy2G4okhkyJW2N7sRA8nzEc5GjxR7DLD3nVe3D/BBvGlJVOeQUBm
q4WKrfR3KxI8ZUm9KG66e9kkJp5xqqfD6RA2MSLYCNhSUbkYTFpir7MbeQfimbXh
LDFXPzW+5EVBrlQ353nHR/Jz5nDr0v01Fw6DAmqPeP2kh0TuOBI0OIWFzkEXfzhv
iXpIDyHYU9LBCXiQOa/rxyxf0SUeCaNInK1t+gZPcy4C1CEPOcVB57otQQNW4/Sl
ND9ThkqvkreZ4GgQzENWgZdtiIImHBKxxcFvbtADdmZ2dBTNgOnXUnb+5lYPYxI2
qjrsiiW5sy5L8X+yayuIkc2soT0I6hk0cjAFhh/Uofk=
`pragma protect end_protected
