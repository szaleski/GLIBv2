// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:51 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
pcCM2KQR2j6Qa7yPTQjo9iC9I7esYwqPD8Swb0/YUft9CG4e76I/RPOP2jFTeFMI
QisSsnBHt6Nb8sfcEL5zuCD81pasfd7knNZnkwCfbiZqvIIshdD+V2Te1avBSB45
fS1+SYiPrTnoEXPpUBiPzXP0ahBV1Zv/PpFyTZ6itJ4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 24128)
eVbOqCI95Ij5LeozGy9pZoVas5aFScvokI/PxlbNk+H7ACbzgA4g4F1J6MEzZvnd
HgYJlrY9MUpft0f8qn9utB2461eAQ+HoIGJv+rpb3/WaqynVj0PYTeteiQfvYj2t
qkan5/AIvkqq8ka2/KxoMC3Au87KKxD+WeVgku2+Lu5hZxhgB7PSMkn3IYIEB8aY
72OAbprh8kBvHo3IPqRmcozplqVf8bE+H7ktmI/TvGLRsASFvc7XfwHTMmSx+pdo
6VbSZdKkKN5xTz7mjqD/9BFWMbw0XLTFSgVihzo6XdhOJ3NIIGmhVox7ygRE38bN
brviqo2ph7fTL1/IGR/hAPOBASmYdAnolLBRUnmyrk1NJxgu5INAEZAesHoseCAc
hpj24L2MlW93p569T0dMxWj5mszREllnwSIXivtpNil/mP+Ce2IHhWBvRrmNiA+U
/zrkdzZu8Sr+Inn2BiI2hKdbCAVPvN4Eo4S2qZQkbn3qH7Ju6O82GF/VU85kgEm/
A3VwqcA98DvWgmOSKiiS/ZlZ82CcLrAUnPm3YXPggRpxyqgvFYl2+auj4IBvwnbv
iqnM8Ne9ZgrAVWIV3YvQ7ePyWJdopOKDw9O4DuCup7pgiX5ERY/w99FX8/qi4Pdn
IsxjrkRBkDNuxF0NRA8c328ZtldXOi4JLneCeD8CR7awwaSQwJb1y0HBqkh3iC8s
wThW27tZnpHc3Ao0CktLSLsZ1IyhSP/1OwrSITXV/qKx0sXIiugNSXd8NaSFn4SA
A2gSjfNVxQynYaY4U72eoPYhlbebIzWjBMZQH0u9j59avug3m1S1IdIZF+ByL3Ok
Qi84f4Zwu1miAsskPYMTiVAEUi3SZ7YWvtqkeK1M/7S5O4ZcXhH1dUgtHiH1L2t7
uOIHZ3vhTDCDd906R0PgFd7zlKb8GVmGAnlM8KWbVI00H3RoL2knTDrocA1KWBAm
wyVqO2Ht+/jw4UtBIjV4acJUnspCFPNBVMb9mMdGwNR38MBiZCDqhN0/JcX46eKy
QcrT5cW/YXUpQbI1trJQCkf3T+HBUmb+pKavMmVp2ZlJ/312lKWePXUH3AbhVM8C
uO7mdaqsjTPaouSEfnFV2v6vEGr1wZvBVy2yxz/JvYmHEqV/Dyn3SfLoNU/XBlHB
pK/l2k41N46JrWJ3ZM8TFz2bRoEIwpWHaHtB2bGdKPLuaM2tTnDvCFnDaYFFXOxH
rXRX6HBse6XvN8d/R771HmXqH2fMKdMeAlmQjEigFWzLf8B82iFSBGRmnLY1aEVW
FoSQiSk+gReDN2idxFHU4VrYwP/rbKOrRwxuMWwY356hpqzakTnwuvnACq/WADkS
G3QTwHl3k7IGQol/J2GU35EK7jjeWeXUiVyDOMrEZvmJkkkFs9EKVk8ulCmT0jKQ
21UISCpmPKtd6HX4uJ4SKg81wu9WZDBgZCwV3QRrNl64XEUa1P7RvOa6K8ri6td4
JluZ9iSNoD7b3c/SkWhbMj6aG86296u5NJS6L/MVBvAPaLwQ7obA1FzWG5vQcOT/
CjMX3pwsIsX95RvgDwBWPTZQOhx0GXoPFjfuGuNlGZICyH1Lop9RRAr3q3V2sMQI
LuzUAOPWQuXFksnor+cEb1jhQMasGDXrAB5jDjhDO3rcYvicGQqGCLHhic69VE+2
ImCw9pbnLtkSq9XJKzzI7TUUNP/3sPhQHixA5+rlO0MrlwYWhQ0McsaK6Q8dQjFz
iliArX04y93eaDY0lPCm8WJRPb0DqYNAa0Ck5vlBVLfilJfRCabqDByQ8KH7cW0I
8IM11/sbTCs8avJNet+dJKUbOpUD6PiA0ATPr/EEKnzlj8njnVwZJpmHQwEad8xu
ZksyiQ5JcuWyr7lcWvOFDbDZR9J56ZXRHs4CuO4kiYRsyG3Wwixl5aAHnUJ7h3S8
UyjDAU9JrVf43ndXJpIv49OFfN11e6GAflBHLT9WY+j7iC9vFIcu4DzKFGvTGy6r
MG2nskP2o2xmAiDFe1U7/zSLbZpBrXP2Q7ycIXmpiPu0H7mVgyq5aTfukQJa3+fK
do1gumUMkG+CNTceVcTusJzbmYgaVWzA6mqzmgdcR2S2QqzHCSEdSrI/p5E3dd+m
dAo88IurOcUc3vnX5RWred7m5sVxfbU8wvgQEVZQjFZATng6OBw479syl8SjHQeN
WihDSB5MeFXplJaU1uVE9BWnxekL2GpeoQTCAAlAia+q4XxseZFTG5vS01FIXoGj
6y5ylQFDezXcuVxCCI4ns/jC6sOdxOAaYdlGFeaD4UHdiEyGmJoq5u/MxCsrEswS
Ek3trBUT/soGGqVDRXkOatjwFJs8iP9tHh3+B85tO+Bl4F85wAh4wY+Sk7zyKdpV
yeFfCTNgQ+H1sS1ul4cG4VJEPnJzo/jwp0EFp/YXwh2h77JR1DwPsMJ8mPVjd+be
SZtMHFKLIrN2DCNuYH2bwcWSHP1M3K1RAsF9TEOcuW1toaVySnDI0X4InQMn0odX
M7he5f9wZmEll8S2+8BCYShm06AKaUkGm37c3CwvbKDVe2QSWzPp5ISlDHDnfkgJ
XSB1zYepKVdifnK6jjPEo4L/LgIRk2jhc2XtqpyZRKI+qsCT6Gp5faikjRc1+2OT
t49+s/F+cxSshnff9vibrDRRmgXGqTifZJoQy+ptLzgFILbTs4FlBE7CD3uTskzA
k8XsK9YGeFLMxH1/2a1usRJZpMjJ47epywWcD2Gf9dXdnQQEL8Ns899PrCKS/4Oz
T/zYHyqE+yOQIb0zKIrJ9N+VXYTNnejoO4u/UurHgdp06uXLz5qsgMbQQ88DWW4Y
V0LN5U3Yx5EeEHyq1+10JkH9tRWGsok3ywW38ZgGZ1Oo1icbbHuFKLAbyRMf0mIh
54Imwu+sExemxXpxW1kJv28NtN4LBY8NPnCNITgxCwqNM8Q5W6/tEQk3cGJMQV0X
szCd5IsQitANUiuiuCef4vSsFiP1EAB/NX8Ozro3U06v//sH8uTkzZ3QIkrOt1YG
D8n4J47VHAYwbrpbrTYyx61nw9UDk0MywjPChUxSoRkTQTaAKxZLv8Q8RDGxLIfz
nUNVvitNpgN/dC+PrWPBsz5s/vawqg+mgoKpNSBsGZGIYYxK8kzCQjz5vUc3y393
KG1KDA5JQXDotSYe6Ch7iSWZmjRAMAlDSoHZimdnV4U6EINlCV1FcyJEDRngNv0T
Bi/QlxugYgtY9FupcD28Ovao/iRxlvf8WGEdgBGvRwOZx7loOXlJ/DFObDp0Hk0w
E2p5NxRgMoU77BKl80L09lzzrBlqH+G07VGm6TvZaCrxHxADybZ/iMZ0VHOy1BiR
ZIY5Ehx17Cl7ltS2rlSBkSKfETnTDQ9cqLuQDnFvW9GD/aXxldjLVJ7DVT3m3nt+
DKABFFn8KEhCGF4WFmoAA3eFXlYS2idDJwP5/65xDqenc69AwYMgCmHsdqNXLU2A
7ncuYorpRFHA8WyL/avUFGoF1Kc6gOnuPeRHSQgSu08h5uxcHTuoIGi2L3vHaVrO
r9l7RCqVSf0U314YrMMXVesziTE8zclg7gdgBsVCLpsqS5cn4EM4LlKkTMI4wx79
0QUcUhZUSu3778vEoqqfymUgY2/kjRgFVB20L6W9AMkxFs2PYEstPoFhz6SxlEBR
IjG8GMZjShpRb1mDGwBUaeJw9E9nUOo76GWEl7NrqDhblJcU2pDmKpfBF1Y7xlDM
Z+hteXZdYkjMy/VDkqf77sePoNK2Fyd4DvGdzp9vtS6xaQAnXWHfBG4Rq2Y/bCGF
Svyx8dEU0N0ejaq/SxqXGQmDHvh4z/+3ENQGpYQDLADQmtKMyxhQCWwKwSPYV+5r
X9aakCaTYz8MRHvs0Ba3KwbpkUUtv7hPJYqYu9djNpqZFq3ObIVrzNv3RNJ+wG5I
Bl9+L+hIqgIHxhD5GuvPqpkD7LYGQQAWIN3bjkUHYX9xptNvLyO6Sl7Kskiq/Bmx
b3QisY3380t4YDhBZ9eC+dwL+l5p8sjjy9phijTtetMTXl/HyvJ1uLS0k9Mh9Sjl
bnEEoivPCcvIEd/9AbQGKSDysOrvUMBBdyXE2FKt4MLKqms6N0UelTk2Q2kHhMAZ
0XfRT/7CLaHDlbO5OjTHnPh/ZLUZNXMCmJyOYLIRRaLMLhcsEa4msKHVFzCoBk0o
G4+2ki/rwDDkcfGWaO/dI3+k37muWWJ66JfTxLXniKprje9xkUSyTVkvW26VXWDA
oEGAPaKi2GtNb/dF4UKO4k3ICjmmd0ZK7z1f2ACOF7SeF2eALXscu3aQLtuJpKRk
cMaNPhw+z7HAWseT/jA7dUV2IMsrv1PdhAXSbOezzD3TPhf+HLo58b2+0qxcAMDd
JwNb65eFprJVKemZsQtugIE45WO51JsBEzai6jJpYT1w8OKZx9BqC3UxeRwhZI8U
UflLTNwMs43TuV5wbIbIabwloRzZ+RrQRHREK8w0fC7hVfE3ORd3l6s3roASsGRS
YY7UIAJHTiVWbT7gVXdAMz5YH+UKgI7Dtc2jGTs4QaDEEeTncZfrzpxsXZ2GY+D9
2hTO+8kn/lqpQwHagBU2nHRDgbl1pe4hMT1HDoKFTBZ4xTK8Wq+gYYA6NvCw5pYD
hOU3wFYn6dRZ9cEy2UCJqwr8dyi/hFg0PkSu3iTVKn/dx2GMuA2lwQ5cUJkqWt7M
1myNJ+n/cQ5mNv9sWXjoHNVWe+ZCfQ0R4iIvxPaVgt8o79TfVym7iGyfry0Niw5Q
q8Ngz2chd5YA/8UyN0fVeVQTPqQJrLejd3m1DXeVjqMfXdFoDBX4qKJVNeSFdcnF
XVvG1KjbcNMWm8AqbhcbFNXg97ZOthOThs4kXghXSL1LuxEaPh3GNshZB7EKc7hk
WWFH7A5Flo7fdHl8cfJKNEAbI7iogJf+PVfzPCLFvJJfnlVpyjsN8/HFe8xzFRoF
MVyBHLAWPusFADXJaL0QAZiSOaIIbvBQLWUIfbdEJJXmPhDhGL/hB+PvyYoIEaHp
XKU5R1AiUw6OkLoHcCbttwxYFUNh7LrudzUSRlIvF4f4lbNRcvrnaYP/5jSOmOxC
YindX+7evk7LBbM7OtO/0+b4qX0gZmaqkDCYFG2sbK99baLEt60eIM6xlnCyzMvz
WFhQ7UFuMlN6mhf5QAWdqhW5ncV8twTEw26qxiHYs5lw74VG50iHp7XiUEnoStE9
zIwP9S9MNbkMHd8DmYsVqM0imJjawgEX7cbMlz/F9CXOUJXksg44jc6MLg0F9T4l
d06YdbSMu+sXL71sUV9CP8nmjaPUeAHHnkK3vCr/gBNdRGMAUNEXn8JkoaTewdxB
9A1w+JykcQBE0mG93Zz7ZnnQF18mgLhvkOGs2LrPrmphKhXHE5w4PIXHqHtFESUk
c8A7XxtXJe+PpGj3yn1WGV5sIJwVIiZlrhHju36xPU5k/HcDEV9U6hjk+sw2SmmF
UH6M/MJs/PH2fGhFqB7Wco2Aedih0UKoVs08X54jY2Uqucu9N9XhQSaFmwgCYK2V
C2topGIJxWzVPRcSfYt/thk5OnxDMu02YpnNjQFE+5Pnd4p3uc7UKCpwVE0zdG+I
9HdlO5gN+l2hZOPd9BlG6DFuPuxLP09ehdhXzbVLsnaOD5GumxTxWc4mXdNKffKt
FCE+rT2eiW6JVhW/Tr+pMhYRs8iK3Us57Mq6alzOn92DNRaD4n3EtYqHWjwGfZW2
xUYNpzO10xsCI+48PVZQX7YIokatKTSQkm6zRuMm84EoyMJpBWeaCSAzl4ert90x
XgG4GVorxwHJ6AAeU6WL5um3iWlmCSV7i20pP7SQM1+qksvjRldD150Qs/Q+mS6F
cik+gKGH3wtyKjHDKLzE7R7zKh0GjNvTK5s2oTCGxqvYwRbbLJFi+hVqVILzQg2o
AN0fi1n0BnQENqOnamxWA5ri5xrvvCHv1oLHq5hyjyCCG90mJUc8xwYmig+ucbc3
LudqYEvffO7R3zwXOzlIinSFPaJ6Dd7eME3NfzxUNQDAwAukFcl9iEorRHQHxlLm
W3oKdghYaPRO/kBlUxigTTj/lQIQGsGhX6CHcbrl7ahNUyBsRsW/NlYWO0hzHCMe
aUy/5eou1Fo07AQWlnT3JHjCNyNgiODKtSf8iV6WxmE52TmRgBKFc0MWf4omoODJ
sjkZMmw5irIm+d1280WaKqiyPoB1nBjF+U3bSo6HZIGEv9zsgOMaRbzuy+3HCzVp
wexK9xcfZnpdz+sb1G/UH8ywc4E+QZ8xtje/tjq/YCiyFKRhM3NDCqvKsF5dv1Ua
XLwwpz1v97BO1fNIZgDsj98Njhfy60J/NDcMWGrcVdPsEIHhj340GxrLAnTCXcQE
UQwzwa+aJnKOUUPEwefrqNkEUb+B7C79OTdHo6NW6qmFkCUTRMGib+MyjmjwqUh5
SDmWg6VcBd06hF84iefixBR7OQ5aR0j21JKPwn1dCmN+uWRPZI8KpC7CQx/eLQkC
BwY45lRTS/720gPL84ytRxANiYRVFhxjKpJ8LgIWEfzS/Yl0BnnAhe/q1LKyoiPC
RHVh4lAEndfMWObPibXvkOi+DJpSMi57oLvX5kAhkVA7+fdI38z+rj4poFf35v/U
QVjIzMMwU2YQYOcpzX+1DU9hhbLDvdiitIwKxxnZ8XzON3a2slaho4q/ZjuTN3Vc
Ls/C4tv2ava0vTfpVSIr9QHDjAyesAu6/E0++TrKdw5FbqkO6eFAFdo0ymEUUo0M
7E14d7hrWgVPnhQ0a4EpzeqsYhDCgTT0QZRFYv+F+9GLqLxG/2of93Yp6z0W2qhO
h3X8DRYgH4FK0B/L2mzhYYP89p8CE7Nzkde5HAJQACz7NTLkGw3Hj8YS8zc42WZ9
aYfW+Xc6fNK7d4gRvCVZGgNAHIKGWY+/O9VCx1dwF6IM9FcKDlMlucN7X8ggOIKe
kScUE1fzGpWQ9k5PUIidnOrOdB4/5O28Zzw3sVo/k7VRzamIenKKrcKWNSWtVe5b
S00oTu5uDVOH2r8V4Nx2sJAvxRxFoIvPX+hbL5s/eJr/HMJ9nYpk2O2vzAL1+Gwo
aKLxGN1tnyeo8vfu1PNAvqn6w8JCdRGku3c3Hx/nGTXw+U9XPeoBZsuc2Qxv6+Qu
vioas8Mw69erjhix8N24QZsm7OUUspgdu2SMgYv0Amt/3l6oQk8o/Ek/4ES6AEk2
IxvCU4lHR1jeznY773svKmhOK0yqKC7U0NEnQrKPboF3QYWZ83Rr1HT4sMy26VIT
bxOSKJFI1uyjN1a/QlUo0XPk4/oZxxXDHCEFF7HCW6X4GJXfUtREnry6CSqDcHwr
QEpQQqFt81yLWu1Ub2JakI6OiVLMiJgP97JH9Y7hccI4pDzTG0wj5L+knVQpren7
8JyihKgPmmHYx6zeLvUOHvCf649ejZK6xiNQNBcpfcBk1MvHe+AoFfOfaYpBqLFA
wZN1q088iSGN4dlqT9zzxzwMUqxJsLBgc7KUifOFnK+g4UbP8fay2gZ32mNRyyqj
MlcrX19kJfdXT1mI27ySU02xC98S67LUfVRtKqy2pd6DcHHi/f3903qC/3clJSZI
mtFT8GBoKD/C2NnLECPrMciJozEZRtdMOxKmVLW4brXZ6G7SbQpXM/rGfIJZyo91
pI10tGHGnHTnZbu3VxFDj7DIwAdxYbLWRD+k9rHVHwH4hDSAG8dHsxqkVEKiOe70
yxl6Z1EugwATizUusDFO380QIDJ27usGIhai/d2paYCY8ofsWYR70eCcjffqc8GM
plqsjE9KLqv2TumidxWm1ycFhcwm8z/EoPavr8TB31Lmt5YE7og2guF4oFWUmHku
QoazqZwN0SU3gRKPPAiirEQ45JnQ5sSjfV2+Px65ErLHY7DYdqULbo8tIaWN/2W1
Cebp4+6HBO5aOZ36q6LuTVpEM0Der5hAvvV7kijMES/raumhvVVJsv2J9Cd0vqQ3
Hne7P+CGYO9OYdwTyjSBi4Elb8s0jWTP/3FuE0Rcz/hRxIiAzJoIFsWY5syxIZHl
mBl5a8f3m+VuRSsCReXTnT+dps8WShN7WmqnF4Crysdrc4S/lKHlifEjVs4umHkW
GB5Aw41QQs+5cx73igISPb/PMOCVlx2NCZGGtCU3TCNgy80AVt8nyu8KKJPbK8tL
qL45dFnDNanPy4VHEq2Ow4jU4dGrHL/j1iDPrTJa6uaxBcxH7l8+2C7r9g4A0qE4
O3pxJ+9ouqaM3fY6R5Ch9e7YB5G+VM7Esb0pDb/bVlPbZ9krfl3oCQVFW+cMPtg6
n1ODl11gcTqDZKTbmwgh8HJPNSErXm/Xz7z698yV63c7HukPRfg+KVkkjKf1A65o
zpekQM3CK3Qn5saEd+AkO8cqirr6KYWPG7ywJdXpQSdqi0dNEU47E9fOE87n65dO
3HZ1dyBxYGX17Cn0mzjZvm4Y0z0/ihRns7OTVrerpaWQ7XcZzx+uU6YyrMKw27qc
ltMufOs0awE+w937gqCrxcNQZN1ywFfqfj6e2AINXVhpdiw9k2BM1RsQAWsqz2nR
SPOSAHJbaupt7ZBsQtq6geZOYf8hyBZkWANwln/otv2F89IKC2L/R54RkW/NBAjD
8w7MTT18WZsOTnjKORe11/i/bfgvQ3hts4EKAuvHKKcCz+TlRnxZy/8VapE7ugEx
CYSH/dQ1uB5aM5y1WR2g/n1BHGQmjj0a5tAKGSCkSx7SM2ojnjpagZBsB11FQdDZ
4Echw9L/ts498gBxJc4APmSbEmijn3hol3j8S6qcPkgaRLocU3gvoXQX7xVRT2EU
eZL1AoGKqk3VI95vimHCPrq78BnMfmsaIN+vCTMj7toltsigBxj6UQnJAfnCKSKm
KaMUzT4YGxlUdbcngR3FzawAcAXX+8i868Z91dL/HwGG7jClNau6OENG0ikXpQs1
Spa+G4jY37ecP2EbeH2WkQl73vL8GWIaws+m1VfNBBlBMrrdoL2G4zQ8HH8BEsxT
FRfyM0kUyBstGT7U4BZA1Sx5gQLTYDV2qLJE7XKXZ3yCl/MYVdGbkak5+1nnD5Xz
81VyrmGbA2hFSDYRjdp5z6e5hSjhBrsfXro+I/zVbZs89r7GYa3jt9EA3+sYzRPJ
e0LlDfpNFLHwGL3xQvfB7FUa/yRp+KjKS/RBO0qLADkLo3JHMKloE18+AWfTfdLP
xBa37vtc7LZ9RJQQey383pQcKIS/DgWIj3TMGc4ikcdzGblwb05TeXdOgfv5GlhI
d2FPqqUwHOcW3Uy88TXlmfEYGicjcyVW/AQVafKzl2FxPCttXeS3OB0nFA5kDvtm
L5wMvkN+6nShiz4ZMITtt2rV2sn55jMb/ONf/Sjfrl16baEvPmdRXhLNzDD/sC/Q
z+DQoE9iFkR2bRNBVL9A+WTSq1rUSLdA//MToSkoq751/EGra5bmWVqKKBdlC3lJ
IEa8UqdDJEKHS9nevBOdsImfFfSQdYqogts//JHd5noPwEV3OjzOASY7pupzxsyy
jLH4COt095Oik35aytuvmjPqDJpBEwKzh6OoESg0c/SrOX6qa608Vx5/RFLzYfyN
wh13OXW2imvSun8Dh8DINw8s16x37AiEVITDkqMZGlrR235lTM6C7VD9Q60qhI8C
4RUxc0/Tq4MEC0AOvWEstAPWHbMJUqUOoZ9E6+vzQ53+ThCzAaML3TWwiLoZGF0C
z7HqRvIOI7ijz0pzLQU7D6ygN9K2VxsnyPu7cVHRdFihiHp8HhQXzN235l53NExd
Oki9TZKGd3dJffwVRy6zwsnIJk3FJbhl4XjCBHjovnKAV77vuKgLfN/PUUahSLNm
NV0dG3IXV95Lq6ZaBM/AsXgpwQSQhQnv/KKo4/Xjqg2uU5yRp6h9Z6XoSSMAD3Bg
qp0ZzgvAmuHY6se+CnX1tg3kHJKLcfIhqNdp2BVaI2Z3jMggsRrUsVZqV3JZIQsu
3rz7bxiLgJ7xDRW6mddNbtQ8FFflkz/d+6FsnzBPzKYdMiewuiFP0BZAqgm2+N8A
vEGXpu7JTPaXXz+c7oWK9/mFFzFmsLRQDuep9T0pifBL91MCmBrf5nZjLW1N+v9k
ItTACcO1ekjecjR9mOgPomI6KepzJyTd99Xdq891ZzQ+IDnGQk7B7GgiRvWiJdKg
hv2gKC1cpejq/8TvHwMw9iPBEpInI/yqjfocLEET5atQJEdVs6tIStx6iwrNUFpY
aYzevyD3zYpo0CMQ8cPZcpDPOYLCdlG7DqIlt1xs7vYKfnfUzjhAbRmZDoKkwyZj
l0f60u3scZaxxsxXBKpPu93NDmYf4xJu5bmCg4qFmlIcNvqYJapZktDtsmketp6Z
8ZP9TWJBIUE3991VkDSRSLJDLFFkyru2AqgC1zochsiBa0r8MnaPocEOmym36CR2
P4Mf1VUG1C0ELfkwGDsp8X16AI5ounFPsINPJWLR+WpQJR5sfxeAMNZLH3CkY9Om
GsTHGrYC+CWR6lgRnHVlJdo1wdd3KAgIo4rFcjDvyhjLnM+T2kNKusz+dUOBUn7F
WezHephsRwkvOOy+SnqT+Pw6JXKAaZSTzq4Wbzvgm07v3rHNvvjAKwhZfO5gMg54
UGmENl8R9eTKG3OFOxV0vKMKyTJPtuqx/TWDuM5c/4c+0lSTUrU71I/Lryc+/oU3
1Tz3oJAfFc33gkb2S0x1Y7DLQZ04OpKXp+WZ5Th10Fr1jvhOPZVmNE4UGNLZkwgE
3ilI0ztO/9nXZMxEI1zi3x1hFHdVYz6XzXVpH/4Z2yC/4GKmpGFhbzGLL3Tku7jx
dre2EzMqzYrOcAKwoD4C2v3XJtYSvvsgcQiYEsp7ewiS60KQbjHDQls8kyrrjxPO
Vham0AsfY9zJ9/usfDLkpwFY5Q5e81MHOVpzQ9WqPdkY4iZ9ApVVcqR5R4Mp5eF2
98nVSheMViMw86iw6p97vZv07Q3l3PlSNL3Nh6G1bckAiP1v9KfWFALtYtYdpuVN
5F9n8JeGG+nNxzTYN9l51EQMOXVIezbG01OmN2oc4X3rNFxOahw9fwPYKqdVsR0j
irUorgu2xq1D1+QIkIFACotLsBDj3BMfmwYwiAsXBuop6dhHcr8UQ3HGB7do4XXv
cGvRRMrl9SoJtNa5/MeWTiYFKbWeHC55WO1e5KcWAwuZulDSdUemdUkjVEDwJ6ZA
44+p2+xHev0pTyH4qe/u/i9GZv04UTvh5qTUKe0rNysy/T9O5cLr/aXQ6p8enTEQ
/LILJRnSFzTGGKh3hKCQBykM0nGAeCu68FVhYRxVaJ/GVH23Bgr5YTe2nVEpMngs
peuJ0xsRn0xy9vm3obY5t+GW/ve2weeTNttEFZVKXrJzJ1p3fZdfnhGBdj/lGtki
hYJqoEOE6DxgP8kJ6l6/jxiofEZCr8El0yybxdOS3PO73nKh14FkIEnLjRMWS50t
9bGzcCuavb/biGq/zxc9WZspGlFNyGBXSbFdXWHsmSxss3NA6/L1vvZGLWHYEQG/
WMGapcSa3Py3jMZn6/dPR9wKfArZ1nf4HbMCvJnle2zZ7g4eGBPo8KVwDMcVkXL3
wykLn8PanS5Q5FM+WuX1QucOyzSxoq1uTGU1jYGwH+1gRdU5fkpGLfBV7D31aNVs
QTMsUE7ckRxobFDyzAvZx8ezEH5moUPpio1A3CTMbYoyGu8PdnUBEegv1aUvPNRw
tZ5RZJZuGU2sPUiEft2NTXjfZTA5a0KaLV78gXzvk5GqHXzNGc4lWAidrjg4k8Jo
ZxDSfeKwVUBE2gTyjkIqJRj3obruFPZDA5IgOeroESczMsLhtVkMFhnu4dUdusya
DskdbGiGmHwiGXVtePqD394ysum7vL86LPA4xoTDnOqYttky7XYsd9lGKfq0mJI0
Sxjp4arJyO45emOuh5H6nwnPhQFdu6fG6+k/NwL77MROm8bNI0A4Hn9ooBcQZYkL
+A7/v8kftbyZWbANvwbHE3JyaKedf8bzkqkrDDrChKAOqaPZ4O4XSSEZMbGCeeQD
g2sf/XOuz9RtHC3Mg5EHtAMYSRtw/d+2B6t3qp3sxqyhsvKNJQBiVA1O9WEuiBYo
4hg3C6yh3wNpVyUKU+GdqTsfPUSqStFsMODw6GrE6QXQYUJXsYpKQB58zhYp8Lw4
6KPVD6RJwukeNj0RaF3sZpkOJ9RQ0Vtv4B8Sc6YgseZtleayqKQWOZg9dq+BjZmZ
bUM8t0nbKrAIFyAsVGyV1xdE7NTrdXfzmAwpefnHu/+hhT812k0i9wJlXvBIKCWL
hPvmxGApOHSb6nHBBdJXS59bukmyxhaer5KmHyHW06bZkA/cL1/Kf7pMNpMKq30g
dcifQ5Z/xZSocBYSuyrEJrmO5aOop0sMKt4aVWW5WSEOVXGzKF3GLXoClYcCQgAZ
3FodsluA1+ueA/ITFBzx7w29+HCA8K/4rkzPAazv73hjHn+CkLc3vRx5dAcEo4SB
ae5+M6YVzybFx3YnNfQ6wCxDZyvEm4Vr0T+BxasBvYZmWn7tEEbPbGqJRAiwP4Jd
PPykmgCbzvCPM/Ci1YYUHoxE3hH/mpiS2hKuydc1eQGy9b+Yre2Z+UGCVETCjxF7
xSEFuv9qP9csQoXv/LNBppI7jiSK310xvRHfgQa6Axhbd5TdetpPnLRHq35wtkAs
wDZsiHlhdJquJlO+98vF3ghNLoienA7j9GpHdAjzfBoM4JUxsWDoraJVl0GLHIJt
L0GtiyHUVPgUYX8fN2+Eu+NQhvaU9qSO71xc18LdcfW4B+d1yVppKVSbopbawZ+5
2k5WJlCcbtRkBlFByg8rc9vR54eucHvx3cgXy/fjsLKpwmtEq3INXy92iRIK0hZX
LQ1Ba0gLYw4Amt7J6v+UtpU4bjlmeYeHBB/CSMydcyFI4G7X6xKazHR5xNLRE6AH
2EMSp9IvgFMcL4QRG5DR3rMs2+n2omBlC8nwHLS3paFqq6N36t2boIqjno0+tsQC
mKrfE69FRcIoAX4NgvPQYLgsvClhKQrAfpk+lTkCkm7pSwcfs6Cex6eavrrWOfcs
Rml6BTdbaSDOJJwyF1UYZLuKuczCEt3q/SPaH12akB3R80BmP15WXLAEyaXAG6KO
MYr2B0KoGjX50Au4YEBM29olumVZxB9z3PFZWr42A1qXLm8gk0G99muKFLouCkN/
Ot3yLfhiO/q56Y/inS2Q6JjxTl0twCYxDw12Elj7vtsZOlceWpZW88oLmWFoX9pN
eNgWM9cT8lhW3Ot7jPHhaOCJdmx7hdCY+bGEBA8Z9nt4DjfBoJr4fOja/JlIcity
Pdvuk8vL2Byw+ttLuOzk/xM0fEdLaKrIwMdj5VUy8kH05oxT65QQcDX1Vwmjjt+E
h6xFqnyqazsAo0O+cOaXUN4cvgeymY0ah5VEhEtlAx8zvF+8bCv5Se/mbyPRcJVV
5lNKBc+bXmenYyJSEHXfuxK9xKTdKUdOwTGb/poWyozRMLlxIRXWduLvcPFBb54R
Bq1O3ZVwU5rMzxJRfpNM4dUnOACFAU0lO+5JB0KFmhy8QUCOXWhOdC7CYEwl25Fn
8kDpDAsplBc3xdZEGxpqVNgpA20vCftSCeKgRhO7yhp8NLSLYJft1QGBQ5UoF5NX
+yfFIBOWXOf6qSyoqnNZanLjp1VJKaZb7kP5vckaWEl+qzZBzRJz6pdGgrxAotk/
cmVZaK7ieFpoO6Iw/8ArpU+tUPrYI9amtkkzIAszkQFL3Rl/BuVPxJNNt2pDFAnD
nOQHHYali+VQsK437ReOvDGNc9C9RUrt9gnHnHwyRzIZBDJYjAoq5KXsWY95g3dE
f2YLM/TcOCKy8/TDvyUxFgP5PmVrqvclbLi2KF1e0r+A+86UN51SOgT44U2DQs19
08QzuU8OI3as7Q+i4J1M0eG8hyvdHnHJqfAY5JJYsa5AviOYu26rJ7sKBFYSyIea
xOcrr83kAUT0jyAztyRU2wneCfVC3hx90YMkHfbT3SCpsWBM5phcTDRlyH6i1oav
lXV2/DqN5WB+k2mS76v1PmywXEIXrgMWBUAfh6UK8CANEKisav/7v8qmgiIVm3Bq
MXE5yTOMb8U8cufbv+zjFEn9Ea39WPqGp0LCUBhHpKqS4wM158cHW2nEsbVysoFn
cOfwgl0cQgJcWiYe+1T4Ixr1S8BVHHT+KR2+jgOR9sW4E/p3StjxQPjA0V1Ugx0Q
rkUxndeK1/iXlV9x6tF9TNSCXY/T0T6x4l5xCNRW583cwJdM3KYoGTrgPSvuqaf4
emmE4YzqZg3tKKKcWw1L0VMjG1Q6mb3XcVgerB2CkRGa72WPQEKPLDlYkO6InKH7
ck4QfMJU+RtSlmO6ik41AM70lFszAxeXKN8PfMzShWXVMteNztbeaVnTidTNHWST
1bvU7ZV/sSo+VNZ/R+NTajg43mGFy3qAQNTFLIHYguq7scnloSNJ1tVAAjrEE/Cw
lxLpwoF+KO9zQm75Mt9b7KIVXtEg2xoU5prZS5qUktsDN59E3swxceclkhi6Ju9K
TKUbUycJKIykTCGZXALOH2nddqbtxy+f3VUV2z6SSqMcHE97bxSleaWrsc3hWnC6
WjjTQE/42YznH+Ryc/spqJqJMA/PcdMfmWRWgFlziqQY0O9m/0mM4Db67xQIsQml
gRqELDj3uCmfxLFmRGOcshLKFd+5FQZEabrpcJDiaKAZcdRpIgTuLTs6Z/F1f6i1
jEhWZw/U7Us0lOYF9rSa9fiaFELIvTP2PnhnGUcwH5ct6i9ZsfFGl8IlydqcTF6v
VQufjLMuwQcauGpnlpS7bri/OyZR6pACZR6GQieiNOKVctvAxxS0hWZpAQiK533Y
OTZIZhqm8rDQmbUOGmycKydrB179kEsSrhMOC2sOB7G+ZFzZ42CcO4Sebq6KIhp+
mfRau9deqD927IjkiuMw6OgJgkxTuOk+s8mDn4ReZPLIbPJtbr81gaxjIfTif/Wo
bUCB12KFXFMbhjQJV+zJ9zDov5MTFtkWxeQkazunlGglAK/+w/vKSD5Tl5LTA6WK
AaW6mDRQKTfgLCOs5Z/JSNNDRasjrzzcbxVAThc5AeU9uUpnX9gMewIAzbOmUuqI
LTBlAzAQvYw/g6MXZpLKdIz6cgZYxC7JWcYlMFaF7I5GznS3g3drfG9lsGwg1XBP
c7VR0XGtdvxN+RKILAS3PiCuvyZ3HRwH3mC56EBnpQBiLkx0zkMaezvhYYEkNczy
D5QYE9YTSwPAy4vj+K6NtWrVo5jskkStSVEM6IDr9Z7Qx7pMbGzQTqQFGY5qyLTn
dHis/xujN43rdgzj9FQFCw0B5yNb+Z1RCkO+s6NA85IBfjc8zDKkjAL5COIH12dA
bwLwTca1i5Nxsqk7zLDhkoIBTTQphexg6pTRoP1cUw4j6JhUrQNPo9IuL/XrpkDi
L/KK9qvVqBLgu5YeP5glCl61WbgCm1c2oTGWHHjGhgu8OL/l0KPdXGz0cQdmy7qN
Ld7rmLh7BcoHCWOtwCx+XOu/b6HIqgueHiPsW26auEfacOBKlJ77nZ05flOf/c5i
lybY80wKo7wGcNp65SoyP/if/EMnGDrfJLUoDBSq8fn0k4/TLvD/HPPqeC0OjZhN
UL/inDxVbHFvVV3nVzdrrzpWHShUEXA8HkLZ7R9akiuKJe1juwflVQF/A95SuTAE
jQ8p7qGesCNnTFlfnPJsgrZt+NlgNI+35G7gllJQ5YIyAzmT4Z1pecvVET/t7Sv0
//XWdHja3bod20CKBBAhmufdlgpMKpWNTt6BBJPfaNCDA8lFY5e3AVMfxBGQB9CC
0+EDFjZBrL0WpRx8x6qrIlgNV4hVlNPSzULbSDf/Nb2D4wCEkFkoecXGeORAxHNN
kFbZZes7gposi2o0QlB7r8Kr2kqSpNnzYsxjio+TzO007Xdhq3Y5sZ452xvtgRje
MYwfH65Koo0xAjNOMYfwn1Qy5qUTRAdenl5uEXAXquiDjpjMoa+vo2cUsiS/nRdY
5N7fs6AkOBXY03m25X06zmTRR6I4J2L0Xs0FFFafQggty2B6lI30Up8t8kZJLZ2A
Og3ZfpL/00MjFso+YksMPzT0kOmXBpOvWnXN6WFP10BOVs7/NoupC2Rq4C7Kfant
q/1AHlaSEVKSE/wggi9KBvHG8J4oOfDH41JYuNAGRpJvG7CGBMWXnGj+IeW25rJe
CpUWjNKd1BKs13u3wMl3djCl0QELp0BtvXRhnIQawNcOjDjcRdA2aTelJmsI0Wrh
z18WbzOuLYC0Xz+7OGUyJB+bQhiUvGsPShFHwZt1StNrKtrBSXLciFUlP9jNLpg+
TaYGwCI4Qppcm+3DwZ+TJ7eKh370H3/uhdRW/5p9ZyZ73zR/tdib1es48bB3na7M
kcjUQpfnMLxYMLOCmkCPhXd4HKZ0bGRW9hkpiz/lN2QYgdzb8uF5P+mHYeCUDj+x
IBBeyXueAQgz/cF4nqXTaY4om1vq8MhnKiAoVzQMdA8FnbMrlZuhAcSGd9QAP5cj
Km41sYWT0tEKKDKWpwC4giRD31ZiFOruXDNm8iQXpmPRjsGipHdve311q0i9RnNy
cdy9dDTFIYxOngG3MI+ihXj+kqtqQ/F4OFMEby+0yxvbL7qjNOaJjGGQtuDBe3qH
xK1q+IjTgTrolsq2xBYpWvHWk5tEJJA8UfkaLapnWDppEfUQ9FAsmZhSv+vMDBn6
6FsUUyxwMAX1mmVEu6UMtBsmqYN2sR+2aamkC4c+3j8Xw8bvRS3R+4PlHj62GhXQ
LwlGYo1R/XbVQ4nBug0swsQdPPIR0EzRomuiPPxKB48XwM9Q+NWNUBiykMd9cZnE
Ab77AOKKsTzVVeurxfPiT3GZHKWi+k3Ak7TAuovV6jh3A6UzuEAXlgqwrQJTXvWf
jlSHpkqzPu/+gzQzmavxuHoWQrdxz6l+Fwv8RSSlVnzn4eMpdiE1wFYZUIec2WP7
hL0388+idjNI19v5UgD+vDDkncM6rqhKo2alevIdGf6n+hNlbIVDrejcQ/Sfr1AQ
TH008VhBzo8K0un9Vzx+vurXW/zBLnGrmFPRRUPJS5tl1bFibrOiZk+3K0XCuajl
UZG85LqmjZgaftmhTpRJHtwHUPStk974bUuYhqjOK2VHa2NzJTFBWoNAtdJsgtOA
9gU2sYbIvG46MZ/H9QhAM8q5DK1sxqdXLJJ9Xls4MuaiENBcbxP2GRu0oWW92o6S
sILEG+kpMM9VFX00W5GiZYyiA47F1olDBjZwbdhsdRhnxzYickXuBc6VnoAgxB02
n+GZDGu4j1Kx2hUNVxoWqm+eGfBcFBErRRJlT3GtDPkuAMvVEJsnm8ZWcHWub3uc
KBcn4/vDiPNiMqahXBTwJ4d5XF79B8N9DCBbZF5o+L5fkrS29g/pLRogws1JtEob
AufoKo1RSAfwRl4rxBQHvzpqNF35HgtphHT5FFDFIu9OlNyBc/KaMmTTFNwcU/3N
qEFeku5n3D4XF+3Rz66qS/DdH3JZkl2lBd+swQoa1epTgKaRmj+QsieYCl51E+vU
fxKx+kpqbqRxAxprohFvRQCTLE5dEV6WaTWnn2JiSEIYjouHSzzin/Oj4XV5rXBc
NDiRyoCfNrNtPHpPmhOQU5NB797oPu2mUaKRsx8rWfIALinH1OGjDy+RN0+voPVk
7XZeqWTGOHXbi21YjgPUOVgu4s5HqtNbmgi7nFrLvyRmmGiS4/YjzAwP272ev/9V
kr0m04spdlVVl/S+NMhWM/cL8kNtkzM5A6Fc0XrA87CnM4yg2aWZDJ6XVKQW6uv9
FiTmbF0/3tQoYZtrt4Obfi0BUjjPyoGutipnkV5beO5OKC4tSBbfW7pKaTvj0MhP
DRvjhUrORrjlDEIwVALYzn4LEFxRw8i9RFeiXGr7Eco5IjBWMJDy4d9T9Qh3Shtj
u5hRdc8TbMGjI9a54RCqSuDef+uoDwIZ2uelPuQrbl2pvr6W/02/NdB0StOp+YZj
HBTXDf+gs9telsm38WO+zJzcNfVwQHdYtLBzaJrNnSgnZneE/u2QNpqrSMDlR2ka
Fv66bhitwtzsUY3dMs0pWCxXV89Ytu+GAvxhVQZgnYQ8Hh5zj0hG2g/6eoz0BnGm
0YaWY6xulCxqBhmYCTgydbFiRa4UyCmc6puZaT/Lo6NhbOsk6OQPEWUfOXgq+VDP
YSxIF1LMIZOSlTeNqS7hPAMvIJ44Jdkbix4Z8RkUY9uKWdBoPgwQF69Hez1zHKo9
RHT0jQqXuuahB06NCKywLEBxD/lT27hV4Pevko/ecCDhoD5+MjFzkjwLi5csEIzE
m9k1X81XfZgc3y59KpY3HFJgYf7NrnqB+OA76GifCV7uA/b6w5w+8NKIwSLP3gxy
Ey05zvjNBa8b0tERGXHB4qZ34gBer+a4diYCt9NoicFzm8wxfuQJ2Wom2UE3YJW5
HmqDcPOqGsOUjEMK6jN1B/1b3BobSe9Ry66QDTify6DUWH+cY/4fcjELeFr9V4LB
1q416ZWBXNoEHpaC9EHgKlE/9NYeRip/ZJ7Jpd7/SSum9KuIgxQP95GYzxi8bzj3
bGiScNw7dNSk86CE7mNEZ0wI4nT7KWrBUAEC+NyZzcbLRRDKe+YPubKFeiwB0hE+
YfmavjSaSsvjk2pocWa9ioKE/zQcvYPBoPUe39Ht+yclMx/Ue0d4rbC+VM+A2y8O
pTJ9BhUIjYigp0GhttIqFqwVNOUl33oHNcgCFDdzKLVN8bOZztxRKCKJyRShWM28
ZFp/PTphZJQ7qxErQm/+6kmMgSG25IYlq1sWoxBHgQYHMcY0pIVRvm+n+hs8mGbN
KFKWkpVmRpHq5y1DbjqfVPCswWj7fNzx3/tK1jJ33pFv9z2owGM+OtsFGFoFQCq6
RoRA3hokdoMJbgq6XlfFkol1YNmdy7n3+JzwMfNa1RSUj96YueNX74DUPL/4AeZ3
j7FyfBhM29vklD5y1laXq6oGe7Pl+n+8pG3b+nqNRfuHahn5V0t1K9TqodQd/udY
bPnAgbFpOt1p15NHtzhnla+oN9sbK0T4HEZ0i2UyqW9FFzZoPLdRGoYWa7mtanwt
ma78wP4Mn3hMZM4+GL2FxPUuc8khvIQBzE5k4iHNNJV+9QCgxUBkGfGX14Bb5mdK
9bA0GPrMCbAktcFQewI5kUMdL5Fk4fbqm/5aHiswPZg6x0JiPLUad00x8/hicKjp
fglnGip6coMWFeEDzHgdh+rop6joySgEC54lBNW+T2C039X5DKmAf80Jv7DEltDd
tiKVW1/jbC3IqBKOKl1QvybbBGiN+gSusxFqMuPYS9nclMVIHJZcNWtl9DhZMqLK
YsDYfUtXlH697D3CV5cvUt2NH41JdIAWN782pJXpbYfKYAIYsd7GCfwPZBldGMTZ
YbbEyPMz88C2gegCaxs5HZASv0b1mpVGhLrd1/iKcN6vjsAgED6tD+hf9RNZoId4
IXJguQw3/286wfE4uyl0UnN0aKcrrICoths3DnTAXeIIpA3xQ4gbics8q0a5JP4E
k+cWfN5AgtIDgZ8oOquhNqBmf1kWeME7PJXa8EXNRPNc+gYS2NQ3Fm8vofcBawNW
1hTrmSweczOFGZcQO3TBPD5Ki4s3nj+2QB6rskISYSUquFNAJSZDOswaMX1rzc2x
bUYZnkjBi53vpfMtBNX9Z67K6/tOTyRikE0RDvpHu+WbQYpuaSpFWa8MV/ena6oK
5//dOCZoCQmxcTa8AB5rwRF1CcRTjcI1erode19iSqMOa6D6vGQXznkAK1ySHyzn
nS/D+k61e8/XIslKxXXoTh8zE6PEU+LexQI+7akdEBTVBALKuBwQOrOwuXJwo+2S
/OeetKv3XiZzpu28N28q8LYqA1mturRy4Ld0Rfq5vOl7p0B4XwwTrsvq19sD+uon
sV0e2EslTem9GuSzuHh1lPVrqtg6tCYeZFd0js1G7nnCwZibZlSN9nPyptZLhI2c
uw+mU+p4HZ1Yia6RTxrbK99yH6ojHwxwF2SvF7gdYZ4oKfsLfGrG6Lb66cF8UI1K
2YeZa3MRBMoHV1OxsVItjeLRBw93E5Hhc8bp+t6kxVa8LO2zVNZVSmnhT2cFXeEp
0BgpEtcNsGtkhHGS1qblNOdELVZIiKiMKNcGkY92rurtjKkGrpfvTYjwQy50/Rhn
pm7TU9M1lMYbxZfSMsMJEvdiOJ67EwASIaxA7N/xpSmPX12aEz+gS/Qiy1fO7Zz9
mzOWQznWeSnFth+Hqd19hDypLTlRfWuWnBNr/8Zsof9IydXmGo3dpafXUcFr0ftW
sMHIg7QOKOBCrpC02pp9d0WeCCS7YOHEQJWWW4/rFr8wRjVxKBl/xYST18mvPKh2
Bar6HQWlGbR/nGV3pfoLc2R76e1f+jlhPYcUpyBWoV+X4GksMR3v4v6VU/7+W5jp
UWwqR85VrLAStQ39GIlOy25iEaeHuKEelYfIXtBQcs91yOshq4krdZc1jWAtPri2
QTvY9z07TRSamGS4nlc2C0Ra+4Nojfgpd3viG+YMwcVRCn46H1xlhcD+NZDLgs10
DXAZyAsTwX8VaC/vaItZ44SEpZr/eMoaZIQg24XPDss0r8H6dpdsYjCWUtNSlTEd
zumxr5tFMBaMikGlsLL6r+Xz5BEIfyVfb+JYeYxVjD7wjQhwc1TusxQhququVW/B
5ByzHrybtg8FevxOJuGxI2PbT+7V5wJft627+tHom+PRncukBYvr3bCKHy+QfxtN
GOMbwFD9SwxcSKukbNm9HVzOrfssvMM8K1Ur0yw15yrGkofbjQ3o9IBLByOV/UWw
YMEcMdsXEVNY1gB9vSBKkT8QRppxg9966WmxJmrL0UEdKRga9DOUqLHnGHd8P1KA
6MT00E/N+cZH+HkMQbdhyLlWWUegSPAnZXfMFCrv0hkERB7vjl0DsGQCbyhcibqo
wBI7qoFcNgLgZANDhEg6EnE/2LA0lQhcNf10d0RIm3OgInRTNv5XCvJdlq6ji8vd
efqZhTLOhtT5ZveE7Unp8qdQEQdaGTIlhZ48KdqwOGFUaF3+JKdajryZvLwgZ1f9
vjC6q5M8nCClboypCr8U2GdkFxsC3UPK/sF4Uc3L5xRi4dfnUn3Sz5ZqUsjepmG6
i5OPyntxEX6u0j0ecy8j57jboJIeh/hRxKUXQZyifOxMmLAfmpU8nr5ewg3eNg3C
NSO++UkCMpF/bJSU/0vdzC6n+bnoVE5PaUxS7wPtgfclr9HL/cv+7MWLVR/Qb+UM
azlgukChgxqVUPVHYJPL7+DYWdf95A6sUMoc7iVzIu9nduJag82S38ViVOYg5J9F
At1evc532yQKyiqU6Bvj4lKdONYWkgE3RkbsEJ4DN/MnR8vpiK1k7nci5HORpyXz
9UZSdH6iCApDUdi2tF41f9K8nCMZDKYTcoc0S9cpvL6wD2ETx+DEidj61/Ev+2Iv
CcCVioE2biU/pDPEINgS8NMW84/IxOySReebRPD0bYm+oXvu5ekMAnAWUVlc+i4a
t055UeJhF2XSapOE/5iaoI+cu24XZjUFKmnq4LbnV4BAdsj9UdqxJd3KmJ9V+rz2
LScrzMClDaV/QTlTuvRxQmZF2DZtuW9i/FtOSnAZi1wPLcOkh+G8HGbJvN9aUdUl
qs7piyVV4lLUENN70sJTztebNHjmaFrpNu/40sV+T7Tw3ot9eOgXDu4hm0P3zs5H
la0KuH98QK5N/lCgYDUm9QiRQJvMoNtNbdCkDw7QnJxg+y6JKhgNa5rVcKtQyQMg
H6bnsz7uHoMzUo8IAr406XXMUCM1C4MlHDVfZ6aj50GkLgeSyVzdG5GjcqK6wJQQ
ePlxTZxJq40Nyc+odNfJRPwnGEMsfeowY4gETWXSE7QwPxvJnMPp+BhhaILWKI14
R78UUv62Dlj+N4eZGlj+D5c0DV03PUmusbxzsRD2CakWnkrKqKB9EIfUcgLlAcS2
gS+rYV8U6zMiHHIbw3LWX3xpqjZTJ+4H5SSEIRfrm2EAi4a2gf8MGHZgWKx8As9e
g0Hp5PX2yWjeuUQxrILNEMn+MMFIXhNpFmQCDKCDijkeQ+SdI7XVxm9egXKJ37Fb
Qg+JKkEeFZuQZiU/87qkYsflPSfx5cnZb6Njg5O4QxwSbC8UYG5yn2E2SlkR3r1s
6RH0bbgoSJj2OiEurKjEvZSUfFbYRUTn6D9zEzOy2CkjOJkwyt4V+bJF8J8ddyK+
jRYnugmvuOgMDKmO1N2x9J/jjfdPJ+oSnwJcUeIlEaW+2qdKuNSv8+WjYJmpomiB
MCW8SaeTR72/wak9faKMChDZfEov5HVpvdzA6GB77o4g2Pt9SxFIM5Rpe0lfeOz3
MSH/bVc76WhDK5DFLLiI+ZVBGrvg6E60CUaqSmTY3zw7bz/w21ecUD97UFBxoQ53
ZyRR8L0I16FIxZ3el1RmRz7rXss96vzTx2/l/FfWLi6hlXm94j4tBhyCGdhDqpAE
qiehav1xxbvjaIP1ptRXQ7KexsAzvfi5XE5EmgD0PjTItyuDKb848El21Mo8526/
dIENdqeAhPtPF4M5lk3iHnUJUbqKz2+dhiFIZlp76bvGGruXBoCAktjH9mG4I/Ry
bYpL0LtmoB7KR2kB5+ZHqS2lABtlaRoyAlU12XTIXq3vInn2sx8rly02a5jjwt0O
ZQsl8zDaQyvJ3VwU7aAjedVcLuGvXtLBBOSMSMa9bEaa8kQ86cXTvvjfiUYKT7kL
CxOzNS/o6WtSLYIfscRCUdBPo5ejLlQdk7NjmMBjyDtLTzd0WUfpbmcU5h/k+TM9
1+WGrd2YWSTsVfJZpOhFcxMW7k0pi0NBmX/yAllKDe0wkK8p6b3SEfKdzwxZudGc
NicFBDLx5l5mfAgZO90Pyg32l+rKpx1EHbWMUriMioji6dK/4e94KGYx5XPNuWhh
EFYsupi4tW3oswqzUwQD+r/lEfbo9VaKYetf75FPuhJ8b7MRlLKmL5OYhglgrh7g
MgHt5Euxv+HlKrW1gzlKryNv4Rcnu6lSG/zniu3otJib5BWTwgGTXL05GGETzmx1
IjjE9Q2UGhfIYNxVUDM9RF/hsARYXclkgzLk7IpO3MXMXbQXcdRPetgRnJKlEiOW
1N6sABOW8DS14c/b9t5siVB24dmPnY5DT86rblRShX6UKZx8I2JbdOa9wjSB1502
k4i3IQP2NGxLyRfouq+bqQkGqpuueRPMY0FnvH8M1QScwY7B4M0Mhe5xHvZZRvn0
8wV/QGnU9zRbIfudAKJeU4WCDcOgzxg5zJYVChP5AGIO7LEfEuSkr0y7s6/F7hxv
OM91C3zK1ok2uP8SuWMRIf4Y2YgHYRGxp50QnPksOe7ZMGFjBboWvZNN/aNRHNmP
7nGVUuGQidAb1FO6fD6//AvJAEmP5IhbjHw85/yqU8IbSyRm7GZoc/O6+7fYlfmj
JXnOS0xOMWeKbo1HyYbU0RaSsS504URjDhtkmvGVRRPxIN1uItOUBBy2r1uZo27D
+YsprxKKhZmhl8NBKkl0v62wh4nlBIOWhBrCAEYSGH4S3EUo0YYmwXhmkHANO4Qe
1O50ov7pcVoHdlwRZ4dB87vgLCR3yHSoGIvtKB9oQtSxPvOih9xbc2+VIfcXllEf
F7ZskYAdd1aS1QUW9xEtHT5oosCjpxfp3hyeAlveikpm/pecd1+NPDBlCJGU7zgS
szbpO1uDYkQUFI5WXr6uye6Cc0wmiB+pRQKvs+5968RsUkXyTLm83DMdwAzlUGCG
hj/oSbLfaTDGpEPErjoWIwdm52ubKzs0tq1BNtzsjY+qE0jjT9E+3lg2Kev/9W2T
doBhOQwYLvJEaFEmoSErNQ6F7WfaLf6wC25CCauA06kmk9VjTSUkheajF3aUD2zh
R69sr6T0qtJaDlMWsj6KxYbH55PqR40GEm3X7dI4PtBihjq77VE/BT421C4JTBJ5
ZFMccJzLYRFd8KQTNrTY5kDbTPa8vZb4lXFHAiipDzVhe2ZFScLNENQXG7TPPyqJ
uQCQGrT+d6pcsYU9T7nTnr3KqMhBMNF2walDnUTA6TFiI+hOJ9sHTB+nPyIVC0M8
Q/DaKarQPmJuV8h58fkd339sXGj7EolgAj7DP5EGQU4sUhD2f7M9zwMzowOctzg9
+K8gSVcIqBiTWg1Zhld9FAsdHLpFQ6j5NFRfnbRTgj/RL3yKOdhSs5kvR4Nkq4A3
MTSQJTjrcahj0BPu1soPCRLNVpTLWbRUIrc1l7EPfQtCPbSi3HybNkTAXe5gwOha
a2Uj21qL7GgOvxnLFlKJjYDba5h3MhVrcSBxEzQfcb4YhXFoxlmBS7WX1SK6dH0y
eVcvoomC8jj/x8utFt/x+4mMvi0nk4waGaj5HhoVj3J+0JBAVmiKXywp95Hi4r7n
sb+i/CMJYr3QZqRP5HGY8ndnGDH6GsFE/axaF5/vXWswt+QlY4OvcFrMvMPvLt3R
YEowDhrGTfPhSfx+f6xzo5v0MtVnOu/ch8rANQ8YWSTVyfBvFIUkf9/qmuyQtlP4
8huXt/v8dWPGeibunbfCLhHFzr20aKM3CoyDNmV+hjrQQ9IbmBlMl/MzwvnZBbBh
2tB9xHep+OgfM3pza09oGz6ML6fD8Vsis1sVne8nm6qCqarbSFWmqV9TEiusype9
L/Nx8qb6LIanOtcMyWIlHrfoXef2um8dQSzew+KmCxsTakiHsqID4pVY1I3hqdHK
IIAcV6BeTEHORldWGtir3vyRgkCOTbCWpX3NNd5UJtUNLDCPReUg9Yozp/h55s4r
qowaZLFFY8R8i88WItcDTBVRlV4TMuklxMwy5SEwSizzPzUrQ4FH0AelHJZjaH6l
II0HamUEl9UappRzTA+sMroUwpfVrtTZTaIqCfJ6cV4UULcYZXAE9j96xRZ8pJSr
DznweA0+1jxGwAfM5N86W//ZbHPXwLqfxkQiwZJkQy+0faygFaiuuI3z/72qJAPD
Rb6ztqktHnSHZzh/SQMtdx4K9Gn+WDPuuYkZ5/z1nKzVkQ5SZdvrT4cPktC75PmX
5QuJ7wgW45/JjZyoDbI0RSsk3wPeSpkGFfGlP4ODHlKaosYhfOtN3LvPoz+VEboC
q6Sb+48CGSsa7LxkC4nAQ6StthCbo6BQ9FXRxRsitNOjc3w8Tn6QfO3M2fO7QBHJ
NVhH8Z8kIfcGB07FFffMheEe+sjNlQdfwRS3PKFFYk5fad8LNiGyawjl/cKH8+wA
i2ZhB/c624VVCUR5U197FCYFZTLJsD/MOdlL2jmgD+ZmzL0uc96is1niXm3GIS2D
edVxP1QzhOtfm9WHunv4fAo2YExx79kWK+VpQGbV/GjbUauzarvy/cuvcK3x5/zA
KR3kVXQ+y4fcvnZ0ieTIvW7IL3ypgUSPGJ5+ZFRm3VwnnmC664Fp2FuV2qKcODC4
Bb8/8zQDd9PGzf1SaPcYO6vNpr/eEIElKJd3nf2ZpX0dRhyiHeSIPpB/JdefNXBr
nnKxfN/Sgn3P4hzRelJp+YBfJDGOar6CRD6OMfppgLxxtu6n4yZqw8w3+AVW1GRT
fzMzoCKrVvCi0yoOTrhsaWVkrqhDFVT4RVkpcwYHVCv+zdrbfvE4kgUWhXFYS+QD
k2cO22m2tkRC4NmNklUk7rAbyKFSFEnU8hy8toGoMuA6xeKQSaYUQif4D55qpKAE
UsK/V2rEcQvc5171iZ9turfhzrnjEqD/oW03XTdXJcoYSFeA+la96ERUAXcBS0If
Y+K04wF+1XsbvsZRP367B416uUSJ3gceIfYwroiRjFLqmI7dtbnBkwqVdPRGM6em
QWc5TKW+EqdgCBuuAQH5lvFfU0FY57vG0oiwvhH0TC3lFhy1R/t/f8m1HogF0azN
/CQH+rjFHIY7oK7xiqwpRNzZKD15CBAR5NVhyG5yfuxT4DCUTFZhKs9vewLzmegH
040XFbA804HvQNq+kS3d05MTpJ4qB0QpYiJgkUV0YZYvV2cRgKQ7ECUMeEU4Lbz1
jg6YCyaKBS8V3Kal9FDTw7lIRPJGghdge/GpmAZkT3i7tUAISdMhHkok1cElhXrR
yNWRceZUojQCRAzRGUOfIq6ZonkKMxcnAvjYIObWyHRCk2QLyHiF51qC2KCZWsK0
DUNZfEgG8MkipzQqbp+NxtQVt9/sUBTzwT1MXn4Yw7H76FkWVaN4Qf0h/SPEA6Si
aB4bSDBSo9JV3eInoRQIdmQfDzMq3wddP72vBkiEwltZcLJu5Cz8OHl4K59YUmC8
uLoUw0tWl3J1CCm5e6K6tP/YTbcol8hX7wwHGLwqBVGQ3TuXvGuaquHzT9WElrae
2IKdK5zUXhi15Zp+2lWfUhc7Ay6w4ARsHHm0oENwSHvFfRSOJIWIc1NhBQMvyzgD
nHPFnLoDjJKrnaEoZkmxQ+3tAWBtD51FMr0rrV/88AWjqRcOGyYLQu13dZjYwzCu
RRjwP4ORG0R8KCkEkS6oYCp87kSIcPzRkR3mkiQQ0IYVUkG5rTaP1cXK9csLMwy1
BSD9wXiukvfk2eBtxqA6ynVuhzqiW0hNm3irjVLIZvAJV4xBgpRN6aWWdhm+f8Qk
5FVv2YC85DxGQ2XxYKBCPaJMTS3gQU5ti8jucmvF8cjH6WHOg9tFy/BX6TyH6hOc
MmJw1G8pT+l7jxd0PT2UPp4/jdWsorSSHEnI2FKjWCZeVqNolv/Y/dqxJVUO3+/t
OXEDVx7FlJbtMMACloAXDdpNmeWkDY0zdTi8kNqbCbPaxwmqhvPzvAgW1j7WmZbE
ugDcEY/PxHRL/SLixaxKOA5WL7ga/Dlw8Ix66JsIjzNEwvIn176FRJlFV5iiB8oX
SYMCvGz0jgEu56yrNUvsR1s8jVDGWuIsLFGtcvsfsc/qlB6GHWep3s7WoCmekODc
Aa2dSJvSy1Ang2NIFDCpWyXCUxvbHoQpMIJ3VhWpT6mH9ttYs+zpvJi5dbtANYbz
cVtsGu+xfY8R1u9FLjosnWxVng8nPv5ZUbwUzWixydKtzMsPZ5xKZg3qFXC64Yp7
0TlXWbyoUtboX97KbrkIKmh9v3qdZfXeD3JReuHP9V6gB/1nhURxFJNqvvAgE6vZ
Ud9+RsHy8nVUCftAAgj4hpeYXkE9WWqUMKfhRFIQ0KmfhIn03nCacKlPC54j81k3
Q0GhRRL5WeG0BD2mSLIcfDnUbrLeAasukQDJWvzvx1D9VeQKxlLAEm42GYKhcn9E
huhkdJCeNKyd2ZlMEl3/WkHh3nxyvuXwWPfsUysUeCztgHpU+vzgSdEkob7dAh8o
3unABJdjc0kJeeuXYj0lmsHg8wlngfpZ+BoE75Y7plHHtkoAtWPkmJw+GZgVXvY4
GAmscnqVE05rI6iiRLytqni8oi9HqOGnn1VfYsoacEZ02UQWteXdltfUGntRO4Kt
ZobXTZ4QoJIPoionLbCORM0K588f+rN7VF5+XudYb/VhTc/aTDNCTs5D51Hv3hyk
8gfSw7sx2FUfxF8m1nc6SP+x/dRTQXqk3YSh6H4yyF5XvpP1UXaCixlmIsCyE8hy
6n9HvXQ55Mu4XzfKzsQ0nutFIRhhy3cF9oDC9HWgun6H/gJKN3/NgR0DyIbf0mXw
UPxj4xu34TnJp4LWHLhmlphANefAffSTCiOlM6IGjUQSJGakizRCj2gRVqMWASEW
8XmPIS81DbgecBFwBISojtEu+QYdrl1Mh1c9kjQ5rmHoLUdPkuTvST02MckTGAqK
q2Wg4OFWU/WIIENRujj1+h8A7GxEU/cgvgsoEk25LyUrYFWZWXoKB7DGvoCKbcE9
gXlWEy2VIY7BQRwdqLVALEZKibQZ4kBqU0rkRJGF6AH/IL/Z5bBBCpLdq1s/8Edw
4eHetTi9j7LmYzz5Skme1SYIgwoxUxN5wmjs0xcobtoP/eoeZWLI6uhwJ3/NaVgm
fLG0qL+X233NozUkV2pTBOPk/uzScx3qZ0Drp2kXWS6GoETcyDIO3MuWRS0is0C3
E22PPeefBtzto6XVT36QT2cEGhgZccLyG8OklCSSWPY9UTWTV3TKge+6q9tMBd89
g8Rs3WpfISVIAYzn2jhAUe3O2bBi7lWQ8x03TxPQf/U6bmYERmbL+VeF91cACwfZ
ferji1vLuHJS5vi3BSCI3FHUoaVtCDD95eorJ3GWb+YsRvqr3DC+ojObNp8haHZE
U+aex8v/Cg7uBlHl1frLHZeAONlBqDXJipfxDWVMK1cIds3lt7m2si9FM79lUL1o
F18Fn9KnMHlJWOwA9GG+3DON3KJwj3XeIH5XqoLsuxz6GU6W8HllLbK62cSHUee7
jF7PMKThKglHsxk3l7+Ura41QIZDhUl0wNQ9ywcB0uvHgSPLIPG1SZio/XVPGWDV
iR1MU6j2R8Xr7Lki3Cw7JPlVe5AZMA6R1xNqGQl6Ps/6SIN1O3nxHWkSbUKctIZE
PVYYZiURFpT4+bS8m4H0PeugbVcV/tWRFjyVAceApckfg5Vdcx17UEqZIRgAZmKi
kmFo5YM/2sorgp9s6I724+iRRwzDy+LUs4gPYBkmvrcyd8ldn2HK+qZaMBKhBf4j
D/68xtFXTzejPhzFO2CPAkZ1Zu7yxy9YetKOQyJ611bzTUQ4bhGMgBHX6EYTMeDL
sTHi5a8hXE2qEB2xvpIDhGw0HlPuJt0CZ3HPNG5MOIe8o9J6H7CnwrCZYWnhNEYB
G4uWppjc5sE5RYqRWXNg019y9VkdKrwtM/PJFDGlo/IMEb0fMc1UkSWe9NuoxEWl
B0HoYsZBo1CZfqfOO7Ny2HPjRXQ7zY4DhRzg9LPV5KZjOMPcyNkMF0szPFgJX2Mk
iEMBBmvuvJZ/1t8d7eZSXXCizf/l/q9mUJCQucgBwCCZheWkBiDJ2ml41Ftk2ToK
Lxi96R3++QmfXCQM7/QWQsD4/PfOZjr0Ve8yinZTicfezORX1UgP1I4gwS5+vB/H
bk9xeJ9eYMZM/5Eo2oqeUDtcYZlSN0z5cwhrziDWepS3wiEMqAnunzUAfDdQDa3p
ZRzIcJWzkvAWL7hMd4R4KluivWtjpaQQcSutjMMCCnWc3hplP5CMQxAA/Yr6sIhR
ZUzToGR4rklIgkcmnfhk3sxyUtTn2Jq12oDhIVCCTrGVxmsWAi0WlvqtBfYiAaUQ
pceqYOUzen4LopGT4d4iNi8AZ4f976TfGWkqtbcfVNsgNdv0M3T9iE8z0Rf+laLK
rKv51zyyJkgi6+Pu+HpoAyRoS7hKXuzG+7YQtkLwtVuoICK0G7CxyaWrizAD5P8x
BGJt7uFIWDQh4mLzV6ZaSQ+aSzR661zX6+xMIO8ywhGSNYnExbXT151SsZL9draV
/eC30MU2OIZxt+LWYYQxSZwf6Kat4wPYes/jdm7wQfmazeWhv4Fh1zAdRSyoR3/R
Bv/EhAxhzD7I2/5zCm5zmTsmleExXIaFSRDy8KvCo47PBB8mR3bNtMdrBowuxQ3Y
f6pQaIRmOZ/N7fNSby9kmj4Ot+S0eODc/kFPkt0S17WDMzySZQp1muW20oyv5Blw
AfeTZniCdeIcFiKG93PGk64RpsEhM4cufgiLpAar3imeAqF5YJmZ4SKF9cyAvTdk
D4qQrmzWfAFGlnMxscGHvHtY9XTDptX71UnNB7Xvt3GP57fY8yqKzsDN/RyKOjK9
nXJnXzfk44Bx4O9DvNylfb7K12eMpaZqVmmaDCzG1Jszj1VLwWQ9YGaPxHhc3vTq
avdnYJ0H1Mtnw1+A0JDRKKkez4h7ScpFcVLkxPEjDywUGirVUpuzVCoWErkOV4sS
NyLZqwwJQdUKYkf70Ya4yny999fwBtl/JB+2buqI11SL0PNm03WRRGp8qFWUsF7z
cgLAUWlqtPH/k/I3FH22xnajlyNFuQ5CieCw51zUtVBsG1uhkSw4UR8x/3PVl0W3
4/fQIriYplOYQER59fgaffZZlIEL8RSKNsGt35JYiPdt8CdiIbd16x2HCyBp/dfl
6Ixo3i1aP3+WOSZBkf8uH+PBLu2n6luOqC+TSyLcEwG086ITv56viiSWdh4xy1vI
Fd0gDQRjQave1yPAbJXwYvO+1DDtNoUAFFSpDArEOsgWir9PaiH37Y+LC8Fnt5pG
2rZo6cTNY4G5FTQ4m117UNqIofWtciiL1g1m4Pbxez5w9JCHox7CYymyyjl9Gwad
FHoCCX/zV97s38r2VwvqRHXbANeQOwfc/0lewlnWQIXJkCi6fT5VO6TK6U4MGbda
WVc7leLm9elzYabfQzWnjcbfPwxfP+LSTW457bu7n9YUZF+Y6LnZGm9Q2WtnfcMZ
Kz/iSDcMhdWsQXF+VLcemysE/xZAMgt0hrhPF5ithayyIShFm7q85rQ7/Ev9GJeG
mB5uU8BtCIiCgw/PwJY9GY9fNhKDBY1VE6wIfqiWzEUFg3Yqrz/kL0es90kQiAsH
/vEcVxYqqXIPboRVR0D4QmtNQPDZvgbBflfbgYVXVddyysgEcNcNMOAFBt+LAg09
9dVyKAZbiXq2cVD1U8eJ5fv9tYtKAUaIaclkfW7a8dcoMqsh0jd0jcEsQFwTmVj7
wYzVRZSltPfd0zK2jg2RdCKWE4N3gDdnNqWk8I6YYRZih/qYatOAVd0LEOFHQNaj
7GgLrTSE6tmQIUQBPUwMn9TwmSzUiFnRiPdl8VzEtoSWl0fZfzpAIS9mKt0Cx1HC
lWxw9j+0wGDZw4Xi3Ml+vbE1JZONrCNSdhkdJJjAxPPQKlSum0rLNS2RgS3lhHXd
kVZEXmwEwesHhPiSDiSzy0+7LxA4H1xrrFS5EosgheLY248DFCzlseAeVWYJ5E1O
bkgF/FBfMH5ThBNRZAHodclhvu9cCCGSKWddalKvl6P0GQe80vxwmhXVApj0u5qJ
Ba+ljHeGyObSw1uZKQoZMhmhYvGRV2r66FvulMcpNYo2F5qY1YyomS/79Q3wGgEB
IVxk7rl14pR9ULRmeYg2nq/MCR5ZZkE+BPEjyNVQ0VNvhmFFwoNXOgM4bHzQHW4F
EGTE6r7y9rUAmsR6mKWr/Od+ykmrZuOZGSpkjhE3Pict7qDl6OD0kJTPTiWIOM1e
AkPD6AjTK7kbgscXzdysm8axiRrWa5/1BTvfmq28siQCviIYzGamIkhKnQN8Sr0w
WBLPAdlRRRLXrlKZM2zRESWPfyVWfl2MeIVb/3a/0Wp1BU0FXT5mh10mpz5fA6Bg
c4TAbYdDd23UlWtNTcSs3aKtuuPl1qBh++ep+yCIPws4zixKAXjyWcaXrAPWiQHs
EyJyRS0JFD7M/ZHjwP2Cc3CHpX94OxU+0D37PcQTFrYrjgcRCCLNYSHWcmQLQWow
2bOu/s40e+ZVVao6nfu96ChxIV89ZnYLZ2jwjKNJCnsDFJgtLhFkSLtRrrWLJy93
2ZZnrUdKiyFdGxc5hdEze3/SZGsc+hvJHWYRgj5rkLcQtjcGI45jOiTC8hyQ5phJ
OIywT0aYdWANkHHychOmj0iyKGRFtsCeMpSNra4Ls0naUfHGgEx3hXEoLyyKpLoo
s5wXhAqtd7oQ5yxJ0vtwJBsenc0qM1PvskteOqkk268k16w3o4EGEP+2CgPn/dFM
Obxi8oABLiFfheB0HrEqSPow3HoSkzw2HDgGkh8G6a0+y6zCTFct4ZxuBKUkjvrF
db5lkTB72+KtqlyLj1JyxB6mDUgWJBllSP/grDF0uWhM67QLMt51rLVmq4zv99vt
xsJ3T3Mq2dJbXRkVJvSrT8FaqbmY5gx/y6RtYRlPB0MnWzJbvKC/C4Ja7NLX/Ond
9uloQExWrWWFxpdS2npqvWQcBi1uzwbfa+DqjuC/fSEiTRAImU/2z+bOnuXcgg2N
6djZ1rwC6BQ1FP8gUfEfJn8Ypebzjw6uzafMSvSFCsFdfnq6rJLvecW7yMr+sJ1i
ZtWVhLA3p6QdtDNKAYCRJOBwW8KKM9EK+T+6z7rBmQNJR4b0aW5eJMCMvodwkuKe
Qm6SsWK6ObmDtGTS5vDcvbUGw/JoGKx+9mPfM/736FHvhyQIlqDu3AWX/Ry0UO9j
AmIy1gbesrooavlOuDQFCskEr5+sj7RocyZdXHFwtR0FfBkdgclt/I8kDznbS+XN
sUo8coTXU1u2YWokI7H3puMxssayn/RPlw82/b3azLiFWfFhyJnF5DACC3rIRpHi
LmkjJZwgAk6OuOLb+z8q3ES00AXCS0pwlJMYGQXvx/60ZDU1XQxA361RPq+Y/up9
hImNqTMy7IPWS1okuEcAn1xnEQD2kP68CPQks0DfX78=
`pragma protect end_protected
