// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:43 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
mePWd750NcLSa2j8qZNgZ11DvEDZiPzECAWUadm9mdIS22lIyD5EtAjKoogMIFoj
m4dWPKrY7H5KJYUobYBmzHHFCez3umcsRByEkJ7y3lqPSniwfrj/GRwry7pmeMWl
Ut9n68ZqI1zRrbUXLEyTu89mDq2ngiW8k93jbtyjNbQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 46608)
CDcYMgaJDCeDgZa678Q1GBWIdDP96l3HMDLyVElFfEqLhYo5aw5paUybidrH9O6L
ziI7wtzJ0dTADw/wItRDNb2v+4peSJqJXIiaRUMGwikM+QRFn6+0tW/r5kUfLl88
v4M2mWT1QVTrJQsqSgmCSpUgaCoFoSDwp6b+0S5uQ54g/RsGRrRrOb6ekPs1CqJM
IoLL3WjWI6y6mCyuzYQTiEdcFESfAPOUiIPLb0edh3WTusW4XoJjNh+GkEPsNpHR
f+jvgs3q4x3TjdejP+0h2MjSq02JJkU5Mlss4R0xSOs93UvZfrBpCN1MhF0WyWwu
Art9aZ81VDrACxeGr0SQUWflg5IyTv0WuTKnP1ER9xqbNbLXECccMNFCmOcXHba8
idh25MG5a5kjk+3kQyEg4Kft/ptXNpgfaqTP7Js7uB1STgbJLK6A8RlgYIrWOKxb
9QP6pz2rRJZAmHoOuy7HSf9711qugoDZ6eyhSfaph6lAn64HIQZ/eyyiN93o0ATQ
lwwIg2HLS1U+vexBUHRWD4Th3Xm9rSGupPBPPrDUdla6WZQ843wt3xoGcjsKe3j6
5nVRJxd07iFy8GEuw+RCvhgIRd+VwB7XtaefYQujwfmGaI4A8xtnnGw2X11z5Asj
w0IUjxnAzOFTJSzW5TMMmI+O57Fc0XOm+w/E/t6eRUAdT+lCM5ZWWeSze9Thyi49
f+a/pcNae56krrdfZD6yUEbUDPbxHr/+uvjmEMvOF71/6TsT+5XV7kMBcf+5PvYN
smuJ9elWBEfsJHLjmBrYzUt2BKWmD7e9UUS9e4r0YgkAjBKUWQZVcmhTjqvWxfub
1/K6/PpUmNDr8VzmnoydLip75gP9laG5PG9Km/vrFCga6XWMpDokECLhkAxXWXwL
SJhcVt4o698t8wKmXMBl82UK755i68hG1TQmIeBEQzeoLI5JTTMNuzuI2yzTI9i2
365abBU06yFXPkMOpCogacY0YgA9dNRPhFTdwQpfyWDQOQ4xY16BcxXOPyvZul7r
wl2qdk127mo3JwNotV8cEFRGLuIgYlF1jjaJV/iz/fWFAF+poisY8NVx2+D6JETb
eyEAgMFsD3zm/AxYjcgfENZ6qu4vazEs7o4Qg7J+WimB+Vqj1L8A+jf0ttUhOouU
33wbvqCsIyAIlEGsX6zXmRku7A4ozt3BpAxI4VDYqGnTEzyWP1ziCJU86SkeQPih
37yTEDFQaPp0Mb/BCTDjowIZbW4t/AkISVntkR+vy4jwaQi5u3JQVExEs2THGtGO
YPVkeb/zZ157yjFeFXbYHuy1qLKmwBE0KrIrH8epS53oUFlBHFCTqi2ayft/K0ym
tG+OyuuSZTSMdWNP5NWH+YccX0V0mYZepoPCPA0j5Iavxc1pMsUrxVj4iPVZ+NK7
h9Hu94CONS0hlDjBphtFAmjRBnbEOXJfgMtnUYc1g2SyCMg0lHH1bWLnQwWEaEgK
3DtscW1FnfHnoEiNCXmGLRxEijHO65P3Qkpgd92SMyuzt4Ai5zZgNxlh9lAA8sRT
OLsk+ZPVYU0iEfj4I4MASmSDn/mtOclY/dc26A5hPl1EBjAYxIG+QeeB4XGwwdj3
PQCOmmfwh/Kf+EOtQMWH1XKevPyfLvu7CfGdd26yuZHmcuwsv+AnrYMC0TBPOfE6
1EOwrFvsCbxsc/Qac9EYX9D0DcxYp9TuKz6M0aqvQPsPB8ApU2Ke7XgQqVkOv4TR
Yyug0vm11uuggkbRo7s3RiYSG/GkrT6b/eTkKvq6ZNOuwhdzEEVtOCoGOFP8lkdN
vC6bMZ7yEg2cG1fHUr1kVHzLkmHeZd1mYAjtOTcUtgspeka1joXXN/MD4LLHM041
FjS5XMKUA2BKJsLWThH8wjocrHT79iBD0STlvyVwPo2QseRMLmelLG0T4PaNxezL
dAfM9Pq7k9d4EsbobAWGsTQ0eDywTs8dQsBGoroIax2+2bPCcvFXKYjvQWGNUzdQ
909phdUFdSrYo73IE6PUb4rzz2ebp+I9kV6yXnet27RNoQ5y6MlbAdWddw/55APQ
dFXqNh+4oVk8Ibdxix6cJR3Xsq6vULyHtBJgYOZA4N7USRcNBT1w4PGB8VqNxiEu
djViNy5Vc3ReAFb5GjlJclJStxv6aU3I3JSphYfknVgV5C/NeK0qJjXPkeil3c4p
/RlFbPlQm9I1Ka12TGqNJ3mZtvc8zoCxe9TckX2fWfbZyybvppDrWBCShy9w19cF
N1r5t8wUu7T6/laZj1FAwTgTbplciUrZokVfsIKgtY0fWoxjX6YfC4d7VJ5v61eM
cyP0tiI6nQ6OUKbmqT913yzMriDe8FwHfoE89Dt3jyJMhcWU8yLkIcvp7V+KvuQr
R2noabGPZOz+kGzmJLTtwI4cf/zWuDyAtEvHBu9GeYtovYN+wEdEmIHFZ7E6MJn3
hI1hhILBzgaOPvl7mIChk6bbJRRACq7qTLeZchtjT/hCk5ArXj+u0P1JzJ9uDox0
EzWTGqEo4OjZO1oSnFB19I+8lOHmMuxLkUOS9zZT3T8Bsu1c7LYUa00KlLL1+gSt
J+A9ldRk7hXSCvZ0aV7dV3e0xv/Eua3X9WfEDGjv9exPXPdBkk7enfUWsSSEB10I
PTCntvm4qhtNahVAnU5V05z1K5C0YVg4RSXL/4sXarWzyPjrel+9BXy39OrJ3d/f
sGBcJiGE8infP1qbD4pSk+f61t1tIRuZ/ro3hcGDES1UGnuiMIPZgxZrJqMUI0/P
3+rSkPvF2MlTc84xY+Cqz23zSqzeJlsBxI8xx+2NJY+m9HuDYOaW0hjuX2HyC8Bf
y7fVEiauNVNInjLYrLI6/9VO6xfWskzdYOy0UKgIUFg5An7fOIL2nDOTJdADhmRh
jQp1PoSOdZhbySHdXfIvqdtfl5V2+9OG4ngjO0Rf+VwEvJielNkILbXSFHn626om
SefuprwSLxqTPETKz6WRXPEX6TvAupGqIg8ViY4e4p39Q7JtBDmbMV0Yk0+UoaYu
WoYwfEx1xTmudGSO8oKT/iDBzFXhoRbPH9u12f5CktlxysK6vqMeeK62YhFZ7+gq
UAYizt+480ogMxZM8fTwWjXslo8CXO3binTLXNnM3oigzGu5pJUJXR5LkXSmc81e
Tpc9qG91tt1LDtbPjBr469gGUeSPFXoBM80jIV5FHXs1oRXOfbhxw665YicLFZdk
pEMnE9pyY6NOXXa0Y2GDv05zo7E/ko7mjUJuFK5D76UU4lD8vi6XY6EPrkgdG+1c
G/6tfF1tqt+O4BXXo5KbootyGpjmyztLVPfr/VAxCKC6GThskd0Lfq7L9PwClWG8
HeUAvI3EcBGq9QAP648djR4l17FcE4CFD7D8I14mnfUUOMR0muGMM3CxUimm3yR6
sOK1serTbtKEkV24dZkiSbGjstRsJ06/BGXR0V0HNPsraoNCGvJR15L/YQ7fcqnV
xSzFBFxFSP/dPfwrBuKqPGaT7p3toth1J9ttNCzIiImoGY+rqtseal0BH0U4t1Vb
/e7Pvn84/Qc41gxCAk58s6v6ciIIjGcp51p29+GeynqPjbGcXXuCQ9T+q/0Zdq7G
P/bHJZvrz42+f/ogAgQIuyPc2TUK4a84muLEBeEnHkt5hhCMpSp0J5qnuKXQc5bd
LgFnlATzJoHgQdgdxoC56SQugtPVrEdV07Zwj3q+KMKYzLPNcw15rPVaKzN6Byv7
yXoQ6dFsKU7cIl1YQd0p3jQKMeCdAo6ftzSEIskOD6bHFbt4QnkOlDsTADlhPaBB
4FAT61EUNcmw5qtO+IbUqXl/zbK3MWShRSvMy2ck9c8o5usjMPTBGvR6D35KdJzf
QgwNrzRWwBOfZnwHR505FyDJRXAfVf10KW0LuCTBBrY7Dirz3Zlf7vWfUsVUoAkD
JexiWZab+WiPcFO1Q3FLCWku7X3zBNj6jeKRTKntkQMjvhkmxUqlbngEn+BRLEiX
7yzVldgnLVxDNJcgh7hQPj9Az8ZeQfY3dJlaoiuGPwwEzNgqBZeCNNVdGWOWrIOW
UHGS3u9OvTBel19A+UQBL8WzzUR5mNma35ZUIr9/4PqykAU5p6qtYeJqIXuQy3CN
yFfF7HZyWIqBXXVLtSjL/0en4pJwczq9IEQ4O6AgMJmLxZfuNwqmZUW8ivHaccNo
uujd7N52GGK4fOL+dXnIU5GDF6vY4aKBPbhYRWQr7jI4XudtjrqRuDwh41nmiDD7
Nk08M/paew7FqTsM8AsdY9416YrUAwhlm/p7U878IuMU/YJJ43km4OQMkl+AHKqc
Bxqhy/Uj+YIqWZu635O+b0wGauR+21ItKSe3Ej/gX+HvW/djK5BlwXdULwIUfwx0
UVkZyjZj83ukSPGxzJWkdPVRqX7uMXRp41QnF1Vo7T4hcredZvia6LbCb1iun+yx
EY8NoSra+Gf4W/iUcC8OpkKQTEajVg39iAAJc9N7E/48lnAQ4/i6Mmbh2zXit3QQ
YP72gw24gfsF6DShqH/WXzDfONO53Wnkp1DsaTXrEhh2NjAAXlxPNZm/hxo1s7qy
eTSOLlOmOurflnNdU+YRqzifWGlFha9Yc9ncnKP7fgwbrutj9sLDXjqddubwjPhk
44BmuLc13nQrko1JhXEDcBCT8Rn1YWefwgQRWCoIVu0fDTHa+08CcSZ5w5EpscI2
EfHowfex8xMagixfR5T8nHnmromOcXW5f7Dnp/R9X65uI1ZAitPck+LjlJ1NwnEv
fXWA+6UXECiQ4QIKrrePYv7ijevkSc2v/NoM36KyRJfxyxnS6ffRhq20BucWs5Ol
vJdPnpK0sj2W8Jr95Y4Cl+rtmWd5kF/0VvvfmtP2oNxU7LeZ5s4eEB9MzETOXBFs
XVtAwfJBi74H/64Iz4HuzhWIp0bYwwF3GYuPCVD4RelnVzJbWmVuTYriduPk7MWo
z7HhDYXqC8ShFaCCtzX82RyNVwaO9XppfSEBcKzFpNAg4HBBu2R9Hyyg+gqmHkb+
OlUpvuOlX4Rb1ZBTlQxdaw0CbppMBqjAeLM03P4aFvzgAYq5vAZ+00mehuw5eNv0
Bz/hBtbd6hu8OOoPAlKaImba3op9bcMsmcjT8J7U9pUKvbsiqYlZrBvgIqss/MLc
3TpB9PBHGuck6xYj6YWRY+LpnD7JyyVwl6f21YOcZ4iStRDf+3hPE3jKXiN9Vaxp
GbfXxYBxmAxJ7ucTvwN8ZHjaK2XaKrwYHK7koSK6pUJqTnE52Fqq2/1LZe3o09vj
1hltMjLcU7Kr4tHWhIxSxyc3BNZlsRgfM/JYLuk9B+eykzX8O8bOaK8n0XLR7flA
NKGoa8CnQEOH1VYLFstGg2kOqxi7hfsCPf0dKNgZDwQ9C0coZY/DFI0rGQe2jKvq
qUGrmHNcdaX4QJxKmp9kZyQUvmtGvilvLgJ4MvfHFAcRFX0wm1SzQRwanYukVDsZ
KXj0v1B9KYjlYKyUW2XpVhuSPf6R48feDnNz/KuJTs268q6VET/GzPKIuhkZ3JDo
Z4Zd6kBhoLiP4Nuw5Pk+gdLd6RmVExgtNE8X5SrSm2Pj5HX6641s2Y4igbrWyxvF
CNXGXILOkiiQO2P0raAutuSgLHvZIz84NIb+RdDcLEiDxxz4pxAG6eBzxjHdArao
zThsi9HV/jJBJorgR4VLBvzm8N3WVSaruSO1P1UQvDJJ3APnurg+3ydQ+asMEBu1
rFuO1eWmY7zjfe6nGOlVxtl35YXPBv8bU6kVgR+K9rY+m4P6U9IDMcjnxbKXha3M
3PshehqL+/QTYsZzyyaeeSci3x2GUp+dIvqGF9V5AFIs7fDjsza1EyuMhntS1fjh
3qcbGHPTJou2UnbLdVWXcgIodKB1QxtQd9VxcpHaIXjWf+SeKy6fJp4pIycAVTFG
JuDdzZkIo7bolNuqLVTF8eU+y9mQ7gXwm5cpu52mcGWxV67rPFrFlryutpgGvPQQ
woG1NHDw0I6tUdKkqO/tlgB+XU1+Vd9XGVVS9UfiH2Dszg6FGLNRwqkki9Jd5wTq
DQkHgYQ0/KXFMwGnidgd5AqcBZ2zvwCNmXFS/dJP472lSOdESY0vdh75SlOOI4Xt
kWL3AjMxh3Q/quY6c4veeDaOBitA2B5Xh0RjIgxmpnECstcYR8fYsabo7gYVb1KW
71GCnnDVu8fsR//pvq5pKG3nWc0HtWcIXYvR2c26w//+PQcUkZMWJ5UJfO8t0HzZ
S0vuIizK1pAIxRBDBORijb7/diG+FDDOu7OIIVSzEcpECSXkh6yTTAkWGYPDydm8
eo4Y/4GC7F9d8SPQDsNCcZC5zo3lNJdAxU7Vun+331i71JPRlKXPtZnHquzPn2Q4
ZZXCAVe0W9tD0bBjd90GvCr3hYReS2Zbm8uZF7pTR2UpfqmePuAlsnvZ/7BzMwsG
rpAy4AeIOQqCDm74FCUl3VJ8ko1geM6Ezm1LSP0S5r0KKCLUMNdx45JtiAzt0ahb
C46wlOIZwn1zHZ1TbF7BHRu1ipSahb31CBi8GR2lz/bw8dqYTnz4oNrl5+qTJs0j
b5wyZHuYsfT1X5pCAxakTIMeikWlO5/YEi1g6Oo3JBiUAjoxd03mlvJ6dajyEHbM
1BWEYOtxDk581fHIm8sV+n9QVIehrxpQC1NRF9JFihn2VVP+0qyd+e9zV2q6gYiW
AXIWOg0CLRVjRmsQvSdW80zlbuIRZ6vkfy9+1mXBsseT7Wa32XVy14KvIdFMViV9
vH99g3iQeS+YEOxHB2TGzt5t3NBqPiUEGuW62KuebhCjtuz+yonfS5BiQaaA6RPw
QVpJllPUb2Wgy7dYEIS8VZdHK7SU3lofwQ0Qz8zVE4uC0s9LwwIQaUekpvnLjBza
JmbBZm3xhqcz4dIRgiUhn8HdlAk9oGnA7+BY2DHc9Ypae1hwfh4eHVt3P8joU7QR
6r69t2WC8/y+vJ2/WZ0s1JfPBTZguiUZoiSkTK73HnxphJT2IZDcL1ELlRSPCu+U
KEnu70bpoR77n42zmTpPG39TGFDVPQKMsxbgSWS/yiskYZYza5Vx8ERcuiw3R/L7
56AD24EyJWlMSpsxHnVjQ5thqKD3dcokjFnyRh2RXuPszn4+oCD2iKDdzddDxotI
FH4KLu4EmLGDdmNgaa1/0oU0UrWn7B8AJumAbr6AnUgENPCefHSkp1aGkDpb6ksT
Shsv7pQe/g8D02Xfu56uN/J0emSM/PsIfjOiACfXUI33klPtEwj+GSf/6cC7g/Vf
9sc5437SzGPab6/ZxBRyRBB5cJG0JY5m3oPjto8hMAspeE7+xNp5rP1ORCqDKiUN
4ve2e4NlV94DTBNAyjKIoea6th0L5exNNK2BIYUW4oTJBL+FaRbcRAkiLVZsrVzQ
ZMomRCiavVH5pfsOC7kLkUrVistYS1Q2opHB77poEA637rbXAzG4uH678DckEYhP
Xd0SgZKPGC162GkvDUQ/ElWTfLkLDwcbRAOkDGioD1JZYtYF55HzooeM3s+D4bZD
rLXwg+1235MnexGzNexQWme55f7Rl5JnrVUfrH364G7XRuRowGvbb/jaS3721R+9
yIkkY2F3vGCiLaf1eGEwJJapBIyQgOrupzB4lUMZajgp6ASnqf3qZqMQirOwxEmV
J7ZX5mqYuyaEDsqq4Yyl1kXeJZ4UIsRe6Q3eTkTX5usceX9K/7CJHttVCUcOnR6H
fUK9SHih0hUNHu7PimbO2iDtmCMBEkVN4a8IogbtI0iDao4oC7OHvX/df9XyCL5M
llHMenlrc1XZ7JTpX8yUA2euwqXWalVrJFhwDougsBCVHtquHEilgsRELWixtGOD
p6PkyWAeYSMcgAVhlXNZ6G6rYUxGxf2e0z9wrHV3nJqhXwB2EGV+w1OCkAK3BTxn
Q4FVQu5YE82YWOcZtPX9GXs+sQhSAznn/QWcZpOzCnq9ac5cxapkvItwpy1cfqXQ
pUI+VHtTXhIeekkAzfOR4Tm2Qekp1JoqZZH58eCyV4UGNuSwv2sHwH4i/JisyzHs
zT1xIxbvN8DZpTJIOnrUZ4bSYh/5ubnrAJtyDdcxx2ztucOL+mkQRZB/AWvIAH91
ODKutEo+bEJF/hZBIgiOGFuvBsLp9a01xBjZfy41eeG1fmzpgOsICoZRxQf83wPJ
lZlV9xW7FUqB6hNlntH9GGMSQWhWDsLrSvXVbBW/A3pmj2tu0MCWonZhXRCv7JvR
v6AuEmZTUYBJC6an9avMahEtTw1xrQrMulIxJ9ynl9tWYAMT6KqK+L3I1MAuiHYw
6CKvN8L0Jga6YSaNocRGatybE4pE7Jkr1ORgSbETg0xGBxpoWVC3TZegtdBEtzks
LC9+/fSOrJyk9gCGMnDC8jQ+iTCAa8bjlz2+fkc2GfVN/7DlMvmW3Th65JY6fDCw
Hq2jUjpFhmMOit1s3DVv8WzGNH9o8rZJ+m6EluSCTAzZazkrWhs/BnJuqSYvwv5e
Aa8zweGjh2RLqBeU6iViv7heKVv+3Xkhyyb7cRGMwm2fTvvGR8nqCLhN0xy8PMBE
cPbVhd3qe6wW/dkKssC8WbnnmKivy3q4T5IZRo3yyJLfO1si3TroHpzSSW0zjPUj
VQVkanHaHr53N8M3YFNVX8qwChoyEx0Zur8pUE9pap6L88NJQFhyoWMvGXiZYz57
fQCln1KwDwU7+FrITy0pf6sSJ1IQ8gJlWJ9ehn8WeBFF49i0oZ683BQy1Sr+eAxl
spjTuPDbqg/Q309gVXuwGqSvOIfWHv10ddnMP/0Pcu8VPSM8ju+FYRAVhQwfsU7+
3MaM903D+iNI72wDJoTRuh0u0uAPge96Ddmz90hsvBnPC1cvtFkfGHGGc5OzlAtd
pfEYK8LGynJ81ZABTqs8AW12f4FLemsEQCZBRS2b7EhPBOh8KXwUuS9znCOvewm/
9diBcFh8v9hE5/YTyOq+vufmzYx4GhFss0pWrcimfZWJGIU1JBRBFxUrBqT23bdD
Tyhc5ukGontKvwaM12CrWlQlT1S7AD6vUjljxFsGCYkh8BP4XSWYevafMAd11ZnM
35MbvE1T0IUtuewyfgZ+c90NbAmiEMcXw9QlNZda6M5Bbb2lr1twiO2fFd+Gz087
M9GlMv5ZZ28wueZOtAfJP4C83gk8ugYwTHFQfpUHSXegvTxz6aiVeoEaoiYaQqX9
HIS/PizwahDFXABbbbTOneJ/7S7RonPDdusKMAVBtIumNnPjZYmBqiLVdnj/KnM3
P6e+fjyrzK9i4f3RRI/Gh49xaGwsuJIdN9/lbhzlj+hTkQVP+/yFK7CYgO6r1Csi
/9aAu1hCY3tgC1Nkb3Hb38TBgyHj2or0buKCaZVekfIZmRmsTEUQU16zrVyM/oeB
aqGsiezFLZVMItZo7+BOqqb4A7TOMBGsfi3SZGkVeH7Juexl2PtVpSiwnZbxmFMn
ehE00PNiZm/aTtE6fVjtr9JQ0vqoqtM2r6fhd8pg7VsVFfRBkxCEK2Jf8wY2Xnew
kc6s/h4y8fwDsS9gm7o9ZjG5zkXqRF8SPAnX/BclMAKi82kvCGoFvslI71W4SzHF
1LUcoJ94RkRR2UAvthbZBqH6qpl3pSFig6P8k9unsT49Ui+JlwlkXX8qoiTxY7Fc
SXBHRZvhsfGVEvaY+h5/SGIC1bU7FkW1DmRy9SVKEX1HLBQdMvfKhqOdn5cLGI/S
l7r0xenBs2PoZPocaOpL1eMXECMvhZQLLQ9CCQJBCaMvYQpP91J7+NAT3Jrp7gst
616EpXrinc6/ftSCXrWRHrbb4MTIHvYkZpvtb597xCMhsriujeHMm23iHikWATQp
ghyX/E5nOYCebhLkdUHuBUZV9hlGEt+I3JcxkFKHu/PSHEC6gk92atT660N6xL4m
katlyrN934lCqX82oivQBgqunOFf61VW3/iWjzR6gwEE2DH1tV7Ps1A7OYuxPH4o
ROFkK1a7wZctJEuTHSL+XwQGXTd3fNtyNchVXnQ3FOOV3hZByfm128TuzMeuxRRF
gC8Hpv0VS4oITgPqfD2Mps7Vu67/6UQRl/XhHZ/XM3GQ9KvRfv2N4DNBREqP5I1Y
jgcyIXOpCQ077Xr95MhEOn3E/qYW7VjfE7XfBiZc+lBAp5wpDONg+sbV6gTFKG2v
l8K4X3M9DQ8Vz7gv9F3JPS/QC5RR6dbXPn3YUkrDxcByuZx6g3LVowvQikJeNLSX
XRcyVSI1y7ryiEpZTbw9pkmSt01KWjvALhDxmsq3iaHxv+V0z1VVIuKpV80sBFCt
nTgfLDiEHgYXx0QnMGTqZPSFRU1NS31PZT95jgYwky34eYIzEhu3c4ScjVUgV+fb
Gcbe6IvWsDqadny4r2goDcAXjCSZqjW9KFvmVZkbgUhhTNnlPQKeueG7dXA5pbIz
TByxEELlkLhCIrVrJ+4CGNvx877ndLG6F5GHqahnVBdVdF4jzOeOGo8fwx/mD2Fm
hoqAIM7m2cx6oAAgioynbjvDLbbOZPFJ4gR5yGPsDOCxT65t2vG0a0LIV3iw/RWA
nHdRQXCKJE4fZYvuI7VWdkTU5ALN1jtCiP62Ox6/2S8yg6QeFeqVO/CAGTWiYsyb
q+C/9fLZDY7nW70g56Oo8f+Q6TJVc7tT38yMHUWNsaVO88f5WxFpQV/mcPbLa+u9
ef3AjlzBEotk2eap/SrQpw79Y9rB7Yc8FrtfGezK5vrhMC92seG4cMdUKsn5VZCe
kz1I36FuGtzxx3nkU/r7Cc4RRdoHK9jqAZnVCzRepRvvogCIM14rfB19Oe9CsOQi
RfMazf/q6avz0+G4zvHVeuw2NrG/5jr5fY+W3EVCm7XYZqsuM7C717wdX1f25lpC
DaqgAOaof8mUu5aj4tvULqx9Pfq26Ep3K/pCf7QlROHig7nhhio3NENIKXAFOMFv
i6IV14G8Y3bh44cJprSL40O3WNsTPzE9+eS7QzuQz4BMfh94uhGaudL30vCOmqzG
+rTlem3JhVlDrblyU9RUPK7JvnjGbAIdBMiEO6V2fssjcRsdZwwzW31NPceZvSHH
/ra5NhnYiFlQUU3Rn3Yg/ipqeIO4O/dRhZDDjWe0HgMiH4PcnUqLIh/fgDzch9ZL
9vN/9pdsjwF2Vq5FiVrNdJrVKCFdeN3obLhPq8K26eKacWqXQ1bK57EQG1yMP2hY
Ih6rxHNxa+LMqt4Rx7QDL0qW5Mfnf3UWY7Tgrc1mJrWXv6lTQcoqzR11ZIfoCwcY
t2gvTTor6k6q6hHEl7QQgQC5/4aY+4oLL+3zFkGR2TBB2tpxrSvElD22vusq9XJd
8u774BVO4Ik3rk8T/2xwy+UOOy9LTuHP+orqY3rna+s7Emh1iu2nIAw5xebzpGRd
+3FDlDPaA2AvvBvdxfpoO77SZogCil+pZ1qpzCAZ0bA3rT+FB/zEpdLkTdhEoBxf
c19ChRdTZuiZWnrHGkrSMd7dUQIEC+FkHsXN8Xhc1ZYWPTzqqbgZ4IYuI1TIoMab
3xljHw6vz/401vIxYwjn/SdgBvwpFHl9JUgzhWTpSVUIRcWUTe52FeSf0OojNur2
R2021TbecrzUWpsbiU2f/s6Aerujc43WssmPharadf7eAszbJY5JW+pviLtCAVk6
WuWXKSb8lJ0Rr0VExvCXXV3pjfyV0+MfnyUm80u9INy975o8hO1eXL3Y2rZ6AvI1
3GyN7iGTlvapwLgaNzkddcV4PqSIJ0hEy4cHK6ribcjHKCl/UEQRMakAelS+6m7+
bpb4SBwpDwtbtd3jd6Bwr72jTSLR3yLMBhu3WFcIvhThNxKv9Z0LjQvG79R9sf6h
tHAOYar8sKK0NNS85rxwF+KC6drFBbEK2GNdcMoxuNlp+wZapXB/+Hcj124bzSlO
noOboScwplyRlmuMcWfeNwNiwC2o8w6niSaH8AiLOPMITpOpkqA7xr0BODVG23V+
l1GI2+n+9L6lddK/1nDpX+DzuHylHMsBub2pOFFLlUMNhH+7cFVYPiXdubsScGr+
TeqQD8WRb53MyHRwY2ZUoRVavyWX2Q3L/2JDmOADNjuPLduvqdezvs8dKTQjXf8v
a9KlOURxOk6nHuDQcJzeRmsG/Ubqpeu5E71pH/8a8hwPh4I/3Ux28d/gItrODbn/
chZviWCgG9dMBFYfwpDIgB0D9M4hvDxwCFnFkDgpxk1bZi3BaYB/kjWjnwuVUZaf
p1+/5bYp0SP+XoE50CarpBdiklmRsY+83btgNbfvcEwaRNyLlB8jE/VCMbInEHYM
N5jy6d90GJW8zFVZZ19q+1yBa8VEzr2BX9EpThs9gsncfMpDfQsIJ2TOOyoLCxCY
BhQWam4IbrX5Lvwyi4l1mkfmwKOur32AnGj/Xhjt3iGo9AJPrbQibkQ9207shDuY
AFCk/ulv9Bil6/C8f0dp/wGRYcAtpdBzPKpvXmaA92/1Eh4xmYYSDws/pwhLgJuE
l+qPx4W2oLucAQLPrPXAhud723BlUVf6nL5aRzqKYwWSG9j9gEYYOa2Kd00hHr5o
hgKkbUq5rghb/j9+KG3kFayy+jGb5Kr6aXREPVa0bFI97Wkj2aiYg2dHdH7jv+BU
p71wg9IZxGZxvuq9TPA0YD0S3eRv+8MKv4vk8a/HMP8q9ElEkSppDFi7Ik/EvwH+
hcNf1Kc12fGMu/x+2b+2tgYKAJ5W9ZnZd4xzmeAeTW4jwGWJHu7Css39xwzqrt2U
y/CTGhqJH7ooa47uzmDfC9OH5n3eKIKAfscmT6aDfwVXitIFsUUv+EQmEItfRcm+
aP0KQKnPxSKLFmh248vm4YRTaeiCxii51uWxVxPqowIl3BPHWnjeH9fs+l0O17pH
aHSmBGZYmLAMXgReHzXHhzE4vi6QSdAKfjGOUqcNvgLNAha9f9X+xLspJTNOpwXO
dqSap3UQqSbw+iIY8s9QEpEZILB/7nd0lXTOhC7ReeDOJX3VMIERrKGVIKte0iij
ghTNCFsnCwNd3jtZHW8RLvKyNUsub2xMc/7Hw/G1hjXubyDlZ8L2o58AIVTnnh6m
XAjlo8XcX00SLMljrnNWTYLAGfv81gWUTigRCK7M8mLBb7k+NaMA3kxkbj5J7eLI
XLQdmwoOTyWCVrL4BAoc9xru41vjWNZ9M15HHFm72Zxr9hB9Es4PWKZYuwZfibPI
3Hck4Qo0YywBqBnXPOzSAtLpA4rEOxtiulskuOEbQk/ntI9N10QLoPqkaYqCG+6F
iF9GXY9MHkdfiMgDmnE3h632egE159Ke2tAWiPbU96awb9tzFBjzsqk9k/9dRYwW
iyt8w39UMOLdWrF2+vqCQqkpGslT7q0k+Svkcyn0NXHXDr3vg7M7Q5a4O6VwGtz4
sj5wnRQ05ldpI3JL6oTm3+/Rw0VWAtQZLaFgfUVBASc+EKhzY7y7NX2wbFfWD9oT
2VhpNhMpGR7itZDMEzFc9Lm57A/joWwcfg7JUV2VHyVVCDcuz/QxGwidnBYla2KZ
8TrtnsPUkDf6EI91g+4KPpthw4+DrIepIdvRoExP5oev0B8jfqrpijNDq3gsNgNz
FsEUhbYRfmqpH1dfF5c0dvN2AxVVdv2HHzdxGbkLibMr4eUeaxcSX+VTyntZaVS/
LbyuXeOdRIecUSVoem/WTaRjNCYb1fyvH8wnZrFpfGznMp3Vxs0UFN+2xSs4tpVl
A5mwX5x+wALEijt4wQp0lkgy/oqs2K7RQVSfz812Gzyx4k2aIbz6l8c38cO9mrol
IChuKH1j9y+e9BO7aWNkXliWNyiEWZSk4F6SSWx2MeG8/xXXpqn/8D9PeVzZ+tsn
XlB2bRXwhutfftg31CO3T9oVrxLBaKwJvmnlFT1zf+KgpIm2wVEs+z8Uq49cRqj4
l8oY7Yn1Tt17xsVL74VqJYuig+QYx9/w34Z1kFFjSgmTZ9qOJIOVa/+5e9c9A6+i
vqmtHOwljvG98aHei5WZiDV8xK+QTmduepWG68dKy3+Rn51g0lTCh/DaaD8lFIhQ
ZgjTpYCmKzoAsq6O5XSpzFdNcHJDy5LJ7F2PesSTnnNM6Vaz/eFlza6Ad/gl6X95
iThbfYjw+FxwGI4XySBmVfcoqqmYo7cw3ka+IPD2iy/aKNVbBA2V9UyJPD/X7CHN
oeQdpaoBazv/LaA2Lq6cEp2beAzSrGDE5MgqOHipkumSeRVLcBvPtFkbVIoJRzPC
ikT6esoI0Pnn53GGKIlaCr6+A49VAQwH0r9fq4WJgLdtTUTf68JsXdrd2QRNksqM
oDbR+uRCoWwiU5UrQFGc74kj4C6nYs4Y0GzkS+P2ppW27fMzNhQrpfzt8sTUsQ5e
+DGtqLjY1uPma4Q5L5PYN0WiuN8S20VhT+Qbc0LfS0nyZqC/L5gylSWdptjAwXXq
zvNrSUUc38lBpudV4WxRWDsQSNXZTX2x5239XaUSkIbWW6Tu4bzREYWlkqHLng9w
BDT3tc+vVVFSxS1QER8RuMcntLPwyctYGC4szz7MuVYAHcdpu7ytmOponKjAHnre
dvkAjyeKZdVsv5JbtrADAJ707x34unoerid/DjDC3R43DZXeYBYeLrwS5F7LcuNf
vcRv/UQUfga7uD8OvLJyZGVL1UKSF9uzaSBKe56jc2saplzk+98GQu0NnaVCgYF4
zm1uq2HciIzYxefFNlvD1ROhATCs7AhcjItetWQZmeBqQIHvjr+pRDCC5WLSdlwY
pFFfFt5CjgvkESV8P6qrcz8yrD/EHIHMLyZLBMWwuwot2KPA47CnTj4wo5BBB1tr
r7WSZxbqipu8ppjbTYz7eCTvJeogleq7bve0xGWvmGJhgMgwKwfEPt1nkgzxkeq8
Yl0Z7/Ch3nuUTRGgApDgA8VPB5ueOHH4OvsZhvn898t6reDCBie+9+JmgQBliZKO
3VNfddFLsRWVB/rU70DXT6Nh726twoQSVVnoEgAhLCGV34UcqDBiG8jO5Vs2N1Tc
8tn/E+L5kjFzzpuY15FVYHP7jEyipSxxk0byjMlJ/G1u+TbVlBw4EAVPKQMYzM8M
zTGWbyYvA2ruY651fIdlI2Lezz9bl/9MOfYGsf2OW7wXiQe02MOHLi0MCg1aO0Yn
lBpiTM1q4MFlU9aFmBj7ctYRjH6VBjyfY0gWCxBJVySxsEAker/TVAIFtZNRffHv
WI4Q6Xv0v8zlFaH2tj/58Mxh8Yaa0veNIxTaeKzbQ5FpwK9cT0rBXWmNra9IGLVB
Jdq3qq3NnVVdglcWvvUTcBmqcgWtAOUGGfPzBo1NF2X1DFseBi+tDEh+33lBHMYS
1E/7hBe/gDIxja0e8+jzZR9qAAfVdZDJizfKhvEWCKVWgQPX/b1TVwpbXAShvhps
C37SkEVho8w3OgUKleUwk7v37cn54WBdemIkVqu/QxAiFabgqYJI4XbNAb5BjhFz
PZ73n9Tk3suWvr/I8R/O8406o4i5MmvxzIXyC24SiClKCwk0+NSyi6DZGF/DCVbe
s+PXYs6NB09mjbKzGN86AsQRrxAqaHPyuqzOyy1whwId+oqMCoKpVqFTFYGe1Mk5
/RRV/7zUwedEdJiGTKevmQ2mwCKt+EGgwcJyMcy56bMV+QUsl8uDAetQM6YNxQ8R
rEkW48VaPJda/Ym8Ztz177PkbD0j0+4y7SKIugi44sZN1ZTYGju1Q2n1wH09wXmW
eB1FpAZzs4zX7vUN6oN8JrJsaViK8lPk+uRvCpwYraO0X/yPkftY7x2URBZpzm7w
UFZAw7dyq73Ooheo19bS39iY5wLBBIcoyd0WEA4ZfpXJnatuSGIJ6DE4li22SdDf
KjDhNnqUmK4lASHQGL3VJ25oQySgBiQ1evlI3w7T4zqFumf1p0TlHpPOa7qg5Gib
d1BsNSlUMtPdAFl9Lt1PQ5O9+E7fC8VNmZ9uXvYIYk+2tWnTYv0zLLED/vCBMsqr
8ZoIFFFh6l/4G+E0V/bhLVVkxEmq5oyy0i3QFDNdZLLN2ZNiyDCmF+pQnwY8Gd0y
a7upiRk1ztrks1RFowdqy+ZGGk2Pavuq1HIISbaEeiFPq4jsfFALmDa2gK+yHYdA
ScxmHEmNpJlxUHBu6CpUXRJHL9jSNKh+ttyGaEDlxF37IZ0ejtWr7S23X0NganLM
atD9F+UHf7V//pz5AkYgWRsZ2rPT4yPtZ+m1rkWg4urnRcpRtmUAF2vqMQmLPw0+
1bnDVyr/GoVCX22xVRD84sxHWK13RfZjn4ur8a6GeCtEbH0aaoPFD6WdnYK11CXo
hQBh3fQYS4Pa2AKuKn1QfAANjUg5cZe0WUNhg38RCXq80xa0Av8mzDn9udYlJ03u
7KwuLgE/DoUejEnKnsPMQLwn9q6NmvduWmAcrdmm5ogr7x53QJjxsQlYsKtvijg3
4VTKhjccgkwSwWcx2BheNI2t2QBDSAd8nyGXwbzgeY5/8vHqKntk/64GLxvND/f3
YjFRs4dLQuTUzMMCgpC0KATprLRHR8uemYLok8YjnbA6IJqlVsJWYDMgiulg2J/9
zTLwWDLObwMTpnAZZAA9gEgkrpnhWPMNVoV6aGurv9CtF0ewhx7vtkQMy3W+8OJo
uUjxhaGu0uxhp2B5M4FAiouEz5dE0bcxu771CKzwgHdXEuAatw8ncQq6I6tc802o
Wvc5baHRGIFN5q46Xocicr2CL3jLsIsdUhfD165bZkC2Kwn40jhvdx4uQZezrJQo
JLtx6rjBeFufQfn6ZY2nPodBt4h4lnpL47/ccWgVEpUv7KIVv49UhXQTmREWXcAr
tFhl4EkJYHuXv8dx4aaqPdXigYwhknAtGlbAEktCpjM0mwVXoJAzT41yLhd3yK9o
T+sSsrLymX/lWmPejrbb/DBCmIIKzxJZQNrBZpdAZe4MfVQHsAWJ/89jIIG+vzMH
V/fLBG72bFRnaJYzDlRwbpZ05J+feK6rXqNr5UjC65wqqcK+/1N1yCRsS/FvG+LC
AfS6kx/K7TIrANrP6Aa6+fj6TklsB3ltRjVsjMKqjS2sokCpgdoO+3tLcvOlYOSv
hj5THYjWduLLdWKBr3bfzg+aI3ZXw439wfXRzOIfCIR8xS5jgwVXPEUTQiCXg9xG
qc3MjU8TMTzNjH6m4PnuW7VlSA0NlEZ+dd7ks9QwVNiApokUV8Ex3UTIoQEGgXNo
S/1hPJSt6u39sWMpaXov1nr+Z+VCXca0nCTDw0ezw09JKFhxkiRf1RSRLmpo4QBf
MA+L4TtUAtKhlFj/pP+EDDx6sTucecPXoHLlRby6H4ZQogn4Ty4BITQt1IxBjjE7
rYURTILGJYFPtzk99XF00G0iPRDikoLXgaqIPBNfsATlmBLgybKGQMRwYfbIxE1r
ssEDkcVPqB3jnQlOvD6FTHzY4DLbZRUi5tJ7E8j+nWR69O1r5Tko1vjX7VZKUAsV
M+xhBq6zToYxXF4eMUrAKFX+NneGVLa8rojM8ikKAdQRc+aZckqXVMUVLCnP1FEL
ZwYlYNtTryDGTCVddgtaRG5WN+MG/jfb5ntkiQ6yucAXsI5/lyvRPkNNhNFQJEVs
mqdJXL/ownAegWdHKBEyiANvj1FRYFKaq33tyA8T3LwiEePAaken1wG8TyIGe4KQ
SvhvgU4+Ebz7kK0p+3K795edwFdyXUlgTGSmcAaep3iMKaUVKIXDiLjWmvATPSAa
Mofp7ot7SIZIFTP+FLOp9bsam1qHXhBUvMnudZzU5L1JkGWskaRosiJgbGnqg7rR
12pzPY+nJ3fjTgDo4lcTSgM/vaVEIyWAMERvxIYUWmgAvKeW98Jav+SgWpiQ/gw8
HFX1ogTQeFLw4nkCqyqsphrKe9gRpNfBQbtm0/RKTRX6883trJXVgsbW0Zpu7YiU
AZFmdt4UtKDm2UK6tNmD1Ol4lGYNpWtSmm/N9NYs4cAO1WsuluS9foWVjrc02+zA
S/MZZFBfpO1ZAr83YNUbfyViV2FZ7bbkin6SAJhcyjjzGQaNP0sgxITEFbv97mV1
3JniSHj7bnNxmCEWTOuvwo5LEpMeUkHcxsDJqefdvmwe2OG96sWYiBfYd3pI7WHf
uaIH3pDizlLmuUBuKfyC+Fd54NPe+aJ2fSg74mXMcoMf0mfEkYJrG59YWCC/KFut
VXz5LnbHI5UXUqiZ7mSDfkrLs1ziG3i2OIrhjJo1K2dkSyHzHcnIrDF6BPKCFGnT
C0TZ7cv3pLjZh+ynTFU6O80NGpskOu2cl9e6oWAI2VuhyMfqQbHBpCov+5eDiO+/
9WJTkj/uZIvKTl69Wy1MKLgELQr1J2Pk/PijY0dPqDAUCpDtnZtvp7c4U/t5JEha
ZeL0ZlrGUanbQYiOq2vK/I1CTW8K0K9Y9tMNs5GYpSfMgbE1MmHCOQV2TSut4Bwk
O6sBisIQ+ctix39nXBhyocDYC3siRhbJPj1ps7gzzpNPCOuCybpASaTmgT8EWFzA
OmChHPvI2gVMhZ6/wAP5zJJ7O8KPBdrRV69hgKh1O0Mxl/7PXW+jp9AHBdDEM09t
6vZGqRK0CC4YREmI1vMGVQlNH6+jH5IKHjdFsspAxtP9syo+eXjOWdhzPmHEbafn
M8+ZE9U3IYlhaZIrN/MD/EKkDaCJ1s3PGMKm2d16NOyUxSTqI4RaEzE4gcPRnlsG
ZryGAupPpgPqrcStUXSoL8AIjyeSBZFlfh+Dfm1HCPMbpbyljKMYqdIn2VeHGIBu
zVFNZBw+1HWi5fN08UGgc28m/477osEUQzF2PC3Ib/Sl5WbFRFgCdLxlCaXS1Pwv
QRhwDDX5FUQA6batXO4FNN3zcP7758FfWofW9ZUMr2R9a1lXlQVhSEE4+Bnxoplu
KrPLkLlvV139beoRpQ9UMYEjayRRMpM6Nov30IBDFOJspVj4kZ7drVOhI49RJtTD
ALHl9c3K/E5gx7snVBfYsxjb7DtsHw3LT0XcPXyJpUAh7nrycp9cKJ+0Ln4aBFlP
XbZyL7Y+gqrHjTK717Q32EmH8OHlS8LgcJcxIe5DqBNVKdALpxaWi+n7Bg8BR2Ge
Fjpg+orJ6SpTAARr4CXfbMz4HD8JUm/GyoGO/WzW948wXSfgUuLxzFCZGDyRnfK0
Y5YkdOoofVxQgW0KpdWxPMjNskXZeUwuW5ao6ShdgP2VJQ2aMM33ceAs71jZfhZs
xLQXc/1EkN/HuhcbCVjCNfL4Hf6jBHZiDER5aTdBBxOjF6AhcOEMnqB4KBcMYHxt
L81Y53bmB/sOPSdIchyoYc1Mu3JugPwcR01sGAB+/lD7fe8QnTBaWdFj1P4dVNN1
mpEDlgN2eHGvjPy4UdFT91+U1iDgrb5dqjEL8d0ueC6HdngvXeAMSk8EwKfEYz40
e5LhCMD6hx0gZOzAirGTvU+Nudo/TFms7ZM1Xjus2MgRYo+hIYa2d9GwtZ1IFXWP
DiDHT9eQs5+vhgcT2cgJS+i5m6FVu27P6mx+yZWcd3cCu9xyDveLSHVeaLD1MLiH
hBnr6qL/iM/PWqBKGSwVLWVZl6t5L/adZjrQaF8J4QbMgGLqsGMB5jl+w1cwppgE
I3hvHirAyuIbPNbSVr2G9IfFvqvSdjtmu3MSFBOFw+G52CB2CELhb8H8Hb0GsqGV
X3g4s87VT1PGM5E9U20CUmp7KLAYalrpZX1+L8g9dAq/2zFRa+0Lqi2pScFyZMjZ
dw1tdCYPoGQ/sNVrqugsYxmpQFjvUKRSv/ifuLm2pY9B7OvXmfGazWy0TNqbtWEg
be0tFb9PpI+weYYxrUnIXzbIDnk4MXg9P3V4oWFRj2XyIFu1MGUKAY9gyNHssyuj
W3p2ZeYfWDssgBJWRrqbsaQQCwseMWclykg/AKllxPUAEcmpHJ9Vr1nCFk1BgdYc
dmBLTr0Jom2J8Y8OMw8FAvUtK46cQYcP5uxwr4SuRO1sRY803IS6Qd7QwlEHnAg3
nr6ltBVPDfcfoDBRoqgE1EEJ3ENj/TALlrZrQacCl8GYNgtJlDBxZVJ8YqWkzFhR
Rd4MB1R40/x9dtLjdFIGrUbXskEB2kOnXXkk7Qr6uViN7vaNiZaHnDPEE1aKuUyV
kVnkH8JHmGKbZwzRzhtT0MRqrkL//JZIAVvdCact537Bu//CBGxzpfL9N26py5KI
JMaYteuQN+MXdwFoOErJ2IlxWjau2G24y1zFRySy8qxI3Ey9sVJ/PI5ouSzEzLjx
FCF3VdOOM+Q5qIHL0YCxCuTjjgLBODPqt2/wVEK8yUQZyjiYq3S4o+0eyUhQVywz
cYQpmHz0pdmiwlZHVbGaDOItT7ayzYcLcuogpLDGsPfyZ1Eo1dcUgoTXaLM2QvTU
HvCXFmBoo4Ri/eQ9bTtYq6Rzxul7LibeL+P2IGoWiEQYFTH/RcsCA8mHrNVzo3t2
A71L55gTwmGWZf1oUisFT/TUc5m8X3/eyqM0bojYDA5KfA2sEx6RzJVXC/TagFAF
wg9PzdgxjA8R2lvgGvtbdkWZy4vWw1czAahTMoSSUOaU6821Gsm7PIfP7GMdS26Y
UNMp2JYE/Uzr0cHuYQT1zugO+IeSUoHMVKoxDGczQ8bA0M9+NiPPzPVKxOUNSEwL
uojVWesvBll5akxeInH0/I9cRH613J0lUXazanWnN8lKpWnqa/r5lAfLUEW6Ajxn
h6PDZhtvmW+JQKpQQJP8tlioV9klxfHDa2Sy9MdJ9+7D6aU0tqA9MhDySgW3kjX+
YGgYdkRVyqOpQ8URA5D29dfiQdNqr2YXcQ928DHpVjqEzU95dU9xKv7hZuYeHgFR
2+Vdqzq2cJnnx0bdnCIGpnS3u1jv07GiDUVVyamnOTZWrCoeWYu+keCZvoqnLj1E
p3ntnRtHSiLTR+UnEMGBFZgSOXKXoD08c1e1To/1e0TWNTI/H1rD6KJo2Wwpj0AX
D8RoxcJJvhFd6wGltSDOSoNVGk3NR9UPFnp2dgRN0IZNTei5Tf362Vb2e/Pxyo2A
GbpIn/ae/g3QRIVojjM/FKDqRRwYQCLW+txrpLExSy0Tpxvf6mipyFkkhBIdQEEY
poYs/xl0r3fSwwQpeBlvC1fj0V7RUc12ibEas+xaU6QV/f0G4mUPWzcAz+MHazfh
QPRNbbwHQxxolwY709thwtAKzqhYR3M5L+bH8u92WV3entksCKLRfYHyd/4EHD4t
Tojz0VdoCgvpTADYT0rxZntgsW1am8woJjqbKKWQ9RzFmRFSN4aZoL2jcWFY7Czu
al/CmbD/8S9gbhJvHQfgn0GxMyQzcKsXZA7j2dF158Rpbf4oK54wSJw/Q7SjE1mG
UEtCANrclSldfwtIFMEI36ibx7I/LxFFdmllGbfmlJh0BWRxAOWOqAHiyvcbOTx3
oEnET9NwbeHO4rYABT3UUqPZn9LY3r2cufUBQyd7RFZbiVDYPpcMy+mP23+Sp+Xs
XJ8j9+2sKso9frkdp5lfoJ413XkAZYBP0MWFO1HnHjdoBqa5VSGVVuqECuHyEQUZ
5aJgHzpTEEsJyQK8rb6csrDHXVdaBrpSpNdLSBLnChGqfZ6BBhX8nLHEJxmx+YvT
Z5d3cye68dnSyoSje7BoeKOzA1ImK5dT1PsC6lsXdkdEkqgmjeQv7mTCybDNdk2F
JsCkvoQdq8dk2mMSR98yai3S6ugQd/xc3R2rLziprEcN5+ApWAWmgZY/Dxswqcs3
2R3yoY7BBGmWKeeITE7TonAAbBJSWWlZW8r3rkfl+KvSloBHgoWRHGBW3cpYyAmi
Iedm7p190FPIfIOzgoTFyLLK46s9Xb7g/u6F+Em/QtfJ3n8/GohcIrqQGXnKIYxk
ZwCGYcQB2gBzBvbtdXIWh4miJ1wCLYroW9kKwuUMQhJx8DyjkGTQfXcgDNG+/1fC
LBWrch+w2Yjn0HBSjJmXQvwlcrhYA3duhLe0iX84MSq3i/GkuYPEnFBxHScGRMkz
ZfVbQgLUG5ljIueb7f1cUaAuNqilQq7l23kit+q3WkBd7hzqV5yCGGtvzcQ4F1Hr
vchESTPxlaDmDaKzCOHEiiguXoTAkY/Qz/xhxPxlJOuBqY7CBc45G31ZIvbBtbeM
PE95C82hjOmfGEklYhQikCFYrsufkNtzQEw++zqgMRkbZhJ6y53tE+LGWJgHGxiB
I/EX00myI5SBNESOhITI20yJvIvPQVRMct5RVhou3uxul0pWFWSqvUznRXRoFOZT
yaFSv8caWD1kc/3PLXhqUXnY6/Z36Shj5sLLGWd5hZfHdB3T4zxsaOWOebCnGmZU
J8u01YgwnbMf2ZlVeOrjsWJzBI6BtWszdswqGcxJzGtOFvnMTgCt0/o+tbXj5iyV
rlDYzRfmK9lGv8sSaxVn9B29widDlkJ0yNlMzOBS2LbQYLf5ReuCmYUeuPKZANqC
2zaxkLVG7/J+3cthHCuhdMYHQiqslfbLqrhbRxlWAVGFM6WJ7ryYDWLbUhf8gyjk
Xe7zkLBI69k7nUOo2IvOzMp+vMp2YlNts5JFDVOxAr0PcJKoQoQzQs2rRcld78k+
ne2F6IcICEV+KK0KaKvGBWlmwGnLvkD6slEli1D+PU/EDNGnRFsk310uc8yackDv
qkSJOXn7Ln48Aw4V/20wWnZkO8++gxq6BIQeQaOh+VVTsEdUc3zIOh3gvNjOP2jX
f171tPmrurA0k+Qvl09gWWFNKx2aYWYr+aXR9fhhRvlUgVmfCs9IH75YInL9qSan
YcEbIa84UIAJYHRZ3reLlqAivp4W7UUIpiMoqlksLXlBXBptwBRAehjK5DQHV5Ow
hv0pFH0QlXWp8TP3LS8mUvrsh123TmY3oqypo+ZJbGtfezLoFxHLm5lpRoSoV9EZ
SFV/nVHoYFJ76GIemnTFYhGobb9a4EGJoeXiDw7oDosZ7sY7Dbb0PCDeFZMqM2Kr
TYmdU4veCLv7FGBUrqNW6/vN7nySzoo9dp1d3naMFxLXgrfi/oAekwqoE+1wax+x
ZPp2FApTvdYop0UnuaoV+z3gxeGN9ZYUIiACrAOXK7vkZZchZzv6ZVgOX1RH9m8/
E0JJ9Dd7HmT813XQz01yWG+7ihYZyZnxjNWfDHdya82kPS6UJRnuTjvbrnuFCS1J
hQ1edanib1OWB2pDhawg1XfX40VZEhXOy5mTbFObe6itpm3Jf6psFBOR1FvijA9m
dTKHvfafQm3mffiRWnjMxTTuYv4p8HE9VbjlteSIqin/pEuoslsYRz/1ziGczFVh
xZt3fyUI8IIWDtSJXgM31EKB1v/Pq82Xb3LugoMD9KaL6TLdbXaWh5uqo4TiOtI9
bp0XYcTkcd11toCpolpGjx6MeKMLrqN0JeWufQT4J7qCezcaYRqfCRI8fEFZU+L7
YJBxI4ujgVXg4l3oauRGpxh/wjtsUt3ZaMNxnB6g7sxU7LIHZlAWSrEKKIrxMKl2
jyyCenXF7GFfcaJIVWIjCASiqJ0FyjOEM5SEAiSSrKL4OnUBs1Vt0Ii7oAo8rKZN
lVelstRFEnk4rHBa2J44AstHxchbQ5cBFSz5aBqbk115/2OJWe6frIhsjNMV/j1E
Ap+6Z6kY1geDukwYWvTH88Q7GNYFQfrf/VwdhfXr+TSPeU93qPk73fvtFto7nQrP
yXMqnEOHZbZlDbHJU3XB89wT3PlSXzde3ETzqAaWsmwzfFoCMexaal6HI1RDl5CB
N+96WSmKyBzBGN4Hakcn0UdQMAnG7L7O2kQ7oS3F90gWY/QkPICgaEMi72Ex00QJ
YOpqS73i2VP+2p6mgSlA70KJ3r1PjQUGMon4BGjQd6MPwvQucduGtJB4VE57Mgbt
6kZ2+BbEBNWE/8D0RtJZl2i8Jak5qrqV25OgRkfkV+Xo2IdqEsbSDI+YGdv9Gexx
i4f3dQZLp3Vso0JAsT7l1wcF/ENPT9I9Z9M+kfQzAHS3s5UHN8AOaETtyhx81gut
5YtVnH3xRxs3j+M84dU0lkz6b0WaCP8lIqTXlqfs6Z0AKmPL6viYrvzfYnUDYAei
1Svl3vrwO4LFIcpswzy0Pt3BI29Hjy0tHF0LuHsY0Bl1EDzXle+CpEYX/L+9+2ya
RqWW2sWZq9VvTdUPkRGNikTVsvlubgpULllBY2qT0R4pcvT9cVG9ugiqUtSYYVZ2
cQcEfCGyNZ8abDROJ03tCDUF9g7XQzD7BUI/oMIDEvSJdhZrH5XGFGYzWAog2S+o
Gy9neDA2Z5hLlNH4ZMDZkNmsfzLOl3rcb9bpi6gbbrckqx8v6d4+sTlKl9SjtVA8
/ReFQpeAblWHjIEQhAvdxHDuvhqITJj0L4RtGW6hkSwfuz/QeFN34OBIAUZBzu8W
fxCCXANd4f2TZwDaSfF0tsHFxJVQebpot/mC2SZC70pv35A/4E+J9sUI56LxP5S8
v5pamwG5TR0G2H0dJVzS6Sg+G1JHGxjPT1VGhiz9noP+W/io/P94MsRgL1KS9OWz
VIlS/Y9OTzX6+nFV1CjBU0JScmoihhxhfO+NbU1joWgPhbK1dv99GM7D25vrFm+8
L6/47ZvgDIpvUTHpZVI1sIXTBZ+m792RiuH5Zm/oewv/L5FzD/dkWjsU9yV8/1BH
uAynhLwzp16+LPf+jwI6BAag+TST0KIOhq6XEgj0AEhuNSNwIa4f4UMbUEBcjIWv
aQ2ZLglVHPtcJFEOSI4JqZ4PrSRb2G35uem5ZW5fjl9mhyWtxNyBfiV7r+70QaTW
kzXnAOB4uc5fdhnSXrgQfyiyNCSdYUe7diT93Lra2CVsgt+PVY531TlyKfXPXg8K
PUvCkx0Ce7NkoWC9W7J4kabQ9JGnBnHKGWlJkxjzT500rbC0Dg4WCFOZGU4qt8xH
k2WLvgFWHhv2uEGVo7GPb+5D/YcDWj2juV40vL3YABmDDWnuE90UW7lNSZmkKi7b
Krr+0OWH6/gWBRNN+XDJ9y7XDOAAVXicHzv9cgcNb1/fXyiSa6su1GU/uBmEe6dk
svjBQ7crGh520Z52UFlPYX29GsXXYZDkj5nadJzvKsOFgP+OGikhii9nf5Yir6RL
CpBAzqPLmYo+BtOH7dvVsGqQ/giMOnF+cIGC8wccGrtM9Hv98CyDSTpl7byHUy2H
9nNJ+gE2hFQ7S5ZISX545Ro3DhJ7RzBNf7elHfS+jQjtG0yrWSbLODETj3rbJ3ko
muvYPJg+bXDMb0BDJ064OXFkQZdTNi0jkerhfd3O1D9uhUjz06uoS4K2VTfSM7/W
48B4e8U371hyK4ZtPeSxsvN2q3xwFy++wy5IX5mlzNTkoYwEAJl2oWZXMX0uILAC
OsV9RYJQZRM6QuZs2QDPRx5Bpif8E3o3kt6dpzltP1I5tBp3bhhReNnIY/sqsqmx
jjtl08hvX6ox3By3LjzucC3Omcs3FWhCGBkJ0kTAgomuYTMxa66eev9EO+r2OyA8
5iGNvLbDqsqQJWs+6b6TGgKVgBPXKjjGkK10MYFTx6ulMBv+LiS8NRKo/7nIwZVv
sjkgS48xurrBIB2D8jo7ZZP+nDuXFQZs9hwGWX9hoODp/kZhncwtbEa8ve/oZYOx
bp+lnLsvnDN6sUYEr9hXM8CAHxBGd1+Fx+sNwXKmLq7O44IU1rIwp7g4M85CDrei
C7Rx1NTyLOcXuGC55A+Ecll7s23TJX6W24ULQx/XKmdkgCnu/X7H0HkNnn2ytAZo
KdUVVxaCAhm5IuYv8Tl8kLXNixnhuHVpQQkpraVHoOi0/2ron7LopQJdpNvoUDKV
TlicWq1Tq7B47ki1QsDOXAiKr/G8lC2/w1/14X4REU4PW0YxiCopCzjytRQWbVrD
htpDECQ0uMkx9jlAyCDT5v8MbtrnXlOSZu/wgSGdH8BhRLV22yPx/X1wX4zavGkW
rzU0O4jXOPzPfQr+KYGtNwKtbn/Lng2OrYO0NgNGbDIaV+h4ctjEWWauuH7xlxzJ
Oxu6/GWIPtDMPSpFq+FzPHDcdaG0FRp4W75lFbQKfm1ZMHvbW6YIus87Li9FOmEd
RIS5sj3nvhiphOtbAHdv6sFm5Aqtdkr/yvlAExWnYRur3jNh/WlgD0W4z2Me5GHW
/w258n9Zd6xfi1c+eDOzRQ25OVrnqIxvy8ix6eDGmsTuqxHB/9KMj82uvfPcfMVe
pVtcXTFYTUrT+pHQom6eX6CJENOXpkqurMTV8CqN+Yaz2pZr65uRBz7WGUJfpQUp
SVX8qXHGvZkWUOVLrNWyw0+UHwgfHNtlS9EbRllvGilYVA10dejSGgMFFfuyT/9Y
xL5tvGPU9DZEVicyNniBUF8WuJiusBsn+M4ZDiO9JDsGsO4Y8T0f+dOv3UoWz7Ra
+sp++wx7RCbPfXh/zAkuP51TBqA3g8oNxb0r6tOS5CHTXp8HpBd72RiKowwMMhKO
FA/cyoFVlDYNChDtsFa92Vz3FdT2KpKTZEGgcqRMcw+Mxi+VLimSW6Px04D60MFq
B6Fcr1MM0I0xkKjKiDBzXPmxokX2i/9rhWn1KY6yp7Nz2AyB0dlOjnUSXqSMod8g
Axxy6aOycRNTo6yUirb97Vq54SpkAVk6NaFOby16jhyAdvVSXiWrpEz8jHWfBThR
NKQOvoXbRZy5gq+a+qluuRMiPbzIPOBZC9rpWTt8HBtJuF+fG9NNUmbvWk3xzqMv
8kPlOiKdkG/2vAkgFkJTDvCW0VlorF48XqGIUzGJkFWMfhl3ZS9dGtzdXkix69XD
qLqX5wO0ch2+oVpVdfY9rR5FvdN+4rHA2K9J7AewUQCk1HjxISx6vK7D/u01/Xgr
1+iaiiWCVbmSDUQ9T9fpipcFvXHz+8M9JSoCUqIMUe9mITqrknnhELYCE1Qt98ey
uvvEqKN+HpO7vSyCY/tBjajACUYguUXJdJqzSe6wO+tuA/MnXLJSNWIDL/0MlxsJ
ii6FoSI5sMPeiuza/kmVjDMUXmIQOycSfpt5O2AQqazjyVIKMFxTZC6UPD7ClZi1
K0P2itqkeCrfWofiV6CAKwrVtINAx0AB5hnpgSV61sxFzrTdzVfetjQmJphCNqXA
fBlMHZV48N8ovCeQd4h6jw9HqJcPodK8Tgg0RfzKlHLwir4ijCUxGHZTTXfX2wiU
CNmTaoRiB93b2Evf4+AO5W1djtLij/TbUPVv9vjaUqo+nf470kbvMrU5D3/KQmgS
XDKSNPkEyyesUd+PmayCdtbKR0WKvMPTY/z9JGwMQIATENALL6rcWMoZk7UR2EMa
3s9n0C0o9V/E3ayQD7UnsLACZyj7h6tBZvE1aL4stXdVj/oSRImX2RdEDP1bQumU
3bTBSA0pwjelGU4GtSZo1YlQLginOzMuGr1h1gXjQHOwRu8tfMotwnH0mCdVGNV6
Z9pDHc9FtYP8QSWb7rAnxqb6IygdHN2B4PdrliWLSgGVQh+rGkhhH82cVsMkjMAD
6nx8Wex1x92GVUCY70NhgsdDf2fV85SjG67dolKTGUqEls2zbc/YQhpWvtO3HNU3
xmlOzbZgvXwK1sVzKmFql1SlM0wp5Rgm2R6yHTjLkmooCmcuYnmbAiIcs0FN8Ksp
Nyl2+mukb8E+lMlAYdGK3MDFDTOSd4d9XthWE3YupfripltEhiIKHOnbRbGxGQNc
pXIHZNUhZoAuAkx/8+laQIMhXFIiT8KuYBLz9nifHAHyj+n/U9gSIkPylfjKkPF4
DGflkPX7B6bdfzpV/8m5lKOSHPZK6F+Y7J6YSfTQz7am4YT5T24rUURN+bewSTOL
pXdljHOW1B1wgNg2/s7u6vgbeOXS2kkSwFDI6T1AXNmakaOY5+k7krkJW2WzcU2V
SBXVvWL7Sop36rXrGBJ48p+4pm5O4FTZtfgoRm7Io7Z8ot8RAx1NOzMsvJQ0aOlF
Aer+lhfjTc771T9A6miuOHWKU0vw3PkQ7jCTRBwoghOXbUGlqTgwRogsSfbwlNGA
dM3B1+740hNCKIFKOfAJ/MJHjH8fadVvarVdlyLZLvdRappZ3j4Oog3giV/OhGJt
e78n/1691rqZSRLsZgl/c8Nd07SLVaH3RrGdCcmMgDMlflow86qEUdu7gUF8GefY
IMn+GGfbR46uq1bLIduUSrOa34iSclk8RAFusPsPc30hhYg7Sq/Ad9140TZMYsik
oNTo4TSL5DJhCB7kVCwXKM56SZszXQKTmGY13ju5cpRLBIcu85rzkBjYBmhnlgBh
7wYI7wwQqlP0SbAlGkp+8F2AuFz8fI11KTwMLWsyb+i9vXjJqdj0FL/gDDEsuYiu
dHwWvY3HHQqF+lSEpT8uBx/RFi2uvSEHZccfV0YTEG/JResnn6BcyAuG1rKYPQis
djQdddoj+uibAS7JouaRawN4SiglJpT9NdcQZcrmkxIsbnnFjN5SToS4bZv0rSGi
NXNV5TcM54mdORkp0ix8Mji6gbnGzRHOrAYRxT/LJCKq4eokbN5lBK+I7YDOFPJu
tvuutSK8UZzIMN5DtfONgv+1AtKqcdgshD8eOmRFyiyuNJZCSWHblI3r1emcH5Xm
ZMw/i2LHVRPpWgMXnZq4gm1uFtHUYcF0/zzwtZeYnyLaZsQhhqk1syU18z1n8EeZ
Lt4f0S8ZMX77pSfMWPVNwbb3v2IEut03Sgz3jDwW6ry+4iOR8bofPOjh2ofECb8U
1cWwJRA6AC7USliH74Dc2J5uj0nrcUV8vf1Pp1/NsUdVq7QS2yIM8LNsdMbRfuD7
zJ0mtwdF7LBKfJBq1YPiRBeERPXBUD2UZ2uGrvM5FSy7ATNb2ksAaiBFBYPpe2Wl
bZjdUP81zipRIH3q7jxrbwWHzaYTPvujtbYxJMuGXQGw0vZlhjorO5tCrHcf688E
ZotenXmLUNJ83tpiZGZAPrGNMfXQKK62afVLQkIe4ZHHOzYC1203+MHu0i8kduNZ
RLwPOlD5W0iJ0xdtCVkBgXMDYmiA2DTfLIvd4rAEKh2NNQLh3a2KXjJQtjHEe+CG
8ocUCTUHoBD6uI+o3kuRYaSKU6u9wiLg9fNx0ZS8elKq4OJ23iEvzANUyMdctG/r
H9DjHlmkQI/mPc88ZKakoHk+PExcAsFIJjZ6Haebg8Zc5QAB9nz3d/slDNbqKxl1
npcoa0UjnOJDMJjasMHJI/7Y1kSmh37jDih0O6kWMW+xOWykSJI8Bqzxb11WwNhl
xVeefsR5beClJgToZU+Ol4PKxS4PuFVgzncGJbffZvkPwE/K4CWF+e70UhhUehPD
e6MWUkx4LFzD+1jeZFad7xQoroo7DoZcUK9Lbkd0RdBjrhXLnDw1O/nymYBbXN4h
O7X0QXBhZ7aq0VOFvPOYr8VHFjAAQPl/VjDJcCfgGyxcQYdmfzoUANZkqIgCW+Z5
NTWDWg3OwqafOIma9dSVSYPwN7mI4Jjc5vDPJ5sMtrWmZwLIXJ/bIm7RVv/7RdIE
Zsso8SSmGeMKA3KrPcHzqEqUsgBApF2Au6oZnZzAhEeFyLtTrPQ2XUMaqQ8rzUy/
jfcNAiojSWYUZI8ARi49zpBgwISRqLL4eDI/8SjiUO2JmLFBPPqPaEWBLRyqSZrq
W2yo3LXQD5uO1uSQTQT6Y8a3+myGhnP/bU80mfMy70GGdPW+y7tj6zAK7sCzdwUc
2Ze4FIbizXXl9b6dGsd6A6bIsU/Hw3mSbS5QNJqrj5laWalgz3mjo4re46UZtE32
4cX4h0WeIOQHjMN7reRdZ7n94onEBDnSId1XTNz4iDBv7KzmQOOUDMaZb4TxW6TU
WPxTPDMCWdkmvwYNYopMiIs9B5SPRWAx8kyEmp2o7D298gCKVU/EoUzPUTd5Klt2
urnd6laePH0/VubAyiMZ+b4mp0Yi+JNL2qbNaLvb5E5PVs9E8j5zdO2RVLnxTdWs
VxhdqPrhp+7peGP8lO/zosBUThuyKQqSPtaJlGrMsD6nEe6oU6zIKllzh9WyI1pk
hRzayyWVy0RhpwJarWfMbNO22/PLabghkVUDn3nNsx01z1ZH2FR0/iqN/b0l/uUh
qc+yW9x1fn3WqeaW74wRbsbZdKFDiEDOauZaD3iEEBUaXGRFgaZPITU3CMHAcoVM
kxbckayd/YZvi7PepM7VJ1gyKb3mu2qa0f2oUurYDgXuOG+vjaCy/oBQ/t6FJmwu
mQrZF+1TmEP3MOc7qwUQqUcgk6UzoXQF4uAOzUf7UTtY+Q8wuwbWIPHk3ehqvUbg
fS6+kqw12xqmBzlew/Qt+3zsicjnGHI6TNBRkgP6uxh6MoNpO6b97dP5Q68TRv0e
N2ujCi23/i30hJ5tAPd9r40pmg6Bcpg8XKR1F2s67cZ3uJsbYgD+G2NyZvufS0lJ
eaxQQjyr41fNPyMOQgrTgRQ7suOj/dWvs8cfdJwhL67yvG/PTJcxd+Sh68v7Hgpl
JUTiO+SIWHVYsyHLUJ3j6pOpPcYq5mIc+5E4eM06WZJhYhQUWjDFlcYYfZdesQLq
3Qtxi5URfUCwGlNiYFLdXX9PKo9fCaBc8d3jOBo8TLWfUV0gcDqgrQ4cGkVvWwig
YFLchNxxBsWteHG8mGfjCrAqXBdtBEBVoA5Mdxk7qPrJy9BraXeHBffaza129nrp
KmAgCTmn6aDatWzhkl/eXfue1QPncmxoDWqi8s4SLWc9CLpcLk5HVl/8hnabXCvF
V+t0QZLri+pIWpiGOM/Mf80GN8gpHCKzFHBzAeS+0fuleNeWECQrIRD60FgtQQrv
jgi1/XCeLbS2KvM33ipVLwqTx4Ek/nLNZEav+Nc3Yk7qDQkLKl8Rxr/+fy9pRXxM
x3Z+yGPUMh6qKVBfQB3dVfTo5M1KY5IuILOpVUgqX4+l3yjbe1WV9JH+aS87pNEt
OgvqOdkJifymc5axJCh08H+Rnzl3Az11lmdA4NhDxApjX3VHvd4FsVOpwzVQ2wJq
7O5FkN67edR/HTHC1E1q3ejAQ+YRhDBUkr6avG4+To69YCrdSHOLYarBzWHY51YO
7Z3now63Ooh1zVSVUSxrsYiyrH9dObW9kBNbg0RmkF5c0yWPVozRrblUEM/aB4gJ
kJ5ClC+yziv8vgi+UXHFF2NcdBVU0tXfB81EtdbiP5Vb3sTiByxCMwrRJPt2VxfS
lFSQL02+HUNfpho+WVfR7GesB+Cde33MTZQQ6avj1ZxDmffMoF8EwWWBktt1KOAu
shhrmDWU6mUzVNSkFz9A5EunLn8SQ8/GUcThiwd39RpG8UitcpQcSYOpV3uiteKR
rxNkzzAT9+QCCOFtzef4CgT2nZ/sQ33BjP739Qy6kstdOU9lDpq/Ya2tb3sI91q5
kOrqovoGhT0XxT2MXjcH2OxQfLCpuR3nBhjPkjlTcEL7hy+Gba2VaerYhxKA9ix3
xrqgBc0eJnsxYWI7vuAp/uM3Je+SV6mq9cqpY7QtO4LTLwlK2xflhNReqDpzhVam
TOZXl1g67JV0K27kEUIiYCz43JBb+QEkyMjP8Rl7gcY3h2JK9fobwoY33fDSzgt+
8+FvNMdhEIz2GoO8oj4KoKKta6aS1L65iUL9Ly39rZAtfFDqYEhJ0bIfxkk04Ru2
yS77uB8XQy26RUyVGalGw0FhYLfC71nZ1zlTei2OBXrOw7nKn9dcgMWgFBfTm8L4
jd9r+oXDRgtp9oLS9m2OBtb9rA/Ev7COxF/DYtaRsinbHqGYJj0VpHYo37ZPCamC
pCJ8aU4YbO70bX40ykKMqZksJuukmxL4u5MT5Um70ZbzErBwpf+2bn/PfZbv5uKl
Adp/gqv7tAzhDOgBXGafBqX5K6YjD22k4/FmZukn4FDAHOEiZ8ErhBWLng11HkUI
oISjYIU700ie0zIbTXJkNGbYfDKY7M+/dGsBKM6g9IWPucvzSF/Ve0fdfoubnXJs
vxVjucb/DSsmsO4cxYVkJA0UVG04U69plM9fC+o9QzbDNWdKljkyXiJ+phtYRKLx
5lqxPJkT15LNawa2G5EGnikz2MIIYkaXPzEH0y8F8EvfeYeOTYlW8PLB/u/Yqv+W
hmoPC+dj+3krNjRNebQQd/KwfbxvLAG7Gu9i2X4HmkLMk7oWVOdGE5l7Be27uRUc
2LYnjGimdq+Dwba7CVPr4WeudSMwoL0eL+ZTIWuYpKmcz5Z+OO1nZg8prMfSVZnE
JlVIKOpKAY1B0IoVIgoyNbFfK9JGQXXm/mbYhV/ylf5ozR9i2rHwRjaTJdKKuoDN
OQAf3YCO6+3+ZWDwWGIhwHnCRHkBCOS6GkBHouAUNJ2pC05awCsUZRUBLQfB5rrP
B83fu15tWkbMegAy7912kbZnew71vNjtwJdpS7nruooe12I5OJxk64a/Q7ZZMHpe
SnEycHrnPV1ZaEl2G1X/iuS1hPly1yoAFyqVPoFlmwNJWGXhz9bVZDKrsPBHzhOc
xRo+L3pm/FDTkIKf32JCoTkHflyZtGkvCn3toA5XuztAJU0qnfwyUXbNmN/iLLow
0d7Y0a201PRbXn3WoxXJ2wLjvOPMSoPa//i//TxK2/El8uQ1eGkFD75VcGQ69aqx
OJZKmZx4tATP/SNcR5WxXeQ2oZpvEZThRI1tq3sQGNxHD3YAsSJSkl9pCGzWBvFX
Z+YIMd+ap0JbwH6U167piMl7qI7HM3OkG8gdaNqw0ptRgFBhpx+3l9raBjJOQ0iJ
U9MgaV+PAgTlp8yCtVx8N9yCSz582px9PkyPAfM8t8iVsdSwtxbVYyM+T58Z95sf
w8Ufnh0U1TcWlelaO12KPakl8jV7gfG1OS84xcSHhQukCWTUxSV1mDqVFWlaTclF
2fb7Ub64ZGVDkCgwitKwUwcdbw549/qb9yUX9x4RHGPAbIqjlWiBE02E1S2CFRad
WtyCDBtHTRJreT1ZX2eegPirx9LDJ8fVf9QTF3l5Qr4L5EDW4PvHfjc2Nk4MyBzK
zn0qpsPK51MNOJ3ra6oB8IjeX9WHIPppFCXqoq6PyOneVxOOkB7WsNb2aC4lynga
oDH1lTEYER614B1oa6Ul9x29kXVcQsEiYyLEkFFecIZgq+SvHyT5adkH5fJ5kfcQ
9fPVA+NYNWR36kXxlyUd+dsKFnzHdzx7+R5jD1yufJsutSlo/vJdlyqiq4Rr8JxG
n6TODan2nOTdfgFhltWv+/HptdtJUs1C0yxwRWWBlrjkqOhuhvFA2oaY5SN0kZ3G
D9J1NnPC0b0MqmKBp4Pup557p2qOvVCpOHDi7hEG/5fUkn/n9vBHITiblfv0lZhD
l0PcEsV4iu9PzWW090XL2RacSEQs5+qvD9r+nu6SSqBwJh6Q5vsfIq6R7sOoSGHr
/a4dzJ6bpbfZQLQdldDr8PNt+cTe5fv1SO/q0fk0jy993E3VSAe+9xB7lUoNzWgY
2+k1AWwDYde3j5AUdx0grHOeFhVTrnP0WeLLVwZ+utCUFzZKCnLuokx2ADysQkXG
LznC6xSzfCCV0/68aCmq52MP47nG5mDzbKSFYh+GlgtDGhsp75E4gWhYwmIhwipu
bejy8uhcTj/ZtDGdWebsRqf7TC01KtmFSXozu24zSrkUqhmrML8bBDtn1ORwk2gs
q/W4J/nw8KUFgNHdstUKLK7KKpnAHMFl8Rq7Y9G3FwbeudfvfnC4m07m24u3FYw0
ODzknvnjBvp4HEQSWInMx7nNstAYJY+tooQc/gkaaU+PO8XvZCwp1SvM1jUZlzMD
E73UqKIoviGzxHa4HX4mvP3JHt+k9nkvOWUetEZnBY7OxtQK8yooUgqvSxZPE4uQ
er3KqYfKjQQ6H76c2l0qglFRPfP0sZxB41S0+CN9d+y7wI40QbLBEcQSd/n1Qxog
AQC96Gp51I075RgMO+muByWMnBrpbNLjpbZIgvKxmFjCqXISCZygjDghQuJny2wb
F5RvrcrjfCCOVv/C+fZ+3OrXdz3oKZyZ73Wt+cxLHAc5IqqBPV4WYQcYsuAa6UO2
geFMTcNG6Hkwr3T2/fM6Zg6m9bVeDadB/F2r1kAubawoX2Vk9eaz8Qk/xNnFCcy9
ZA6OpQlKi6N2gXev3gqyfMueAwz5IcqOyrs4OFZ7GR494LJLmboj+ogoAS6+2lDI
uB9tMTzRI3VhLfx8ku8tR5pzzaJaBb4bMA6jlFCfNd5cfPrPeisB18ZfTjMgPPi1
K7uj00OHVtuv//IOaBmFoPF+aCAWOnfc1BZcJl1wljC8EAo0EH9S++c18LbWDTXs
DKYPB/13EDhWArO2nZesRmVA6Wx5ut0/hTOQKC9nj9M5sKlto8PDpGgNx7r7NcRS
IS7gVGF/leznk30eLauko08mnfSgHRLe6oi4efm/DWtXqli9laO+Lab4Fn+Z3s4S
oQJAno+DS6XAdL7QJtxjHNqnPeeSKkV289eqnGcXao8A/9EBi9sUEd+IKqjMHBxP
UsWlfHKLBPFgmSdY8A8QhIICM7w5uYrJ4Z1IowkZv9I/4ZWYi1N0BQKdWTgzDWK2
AVYnc+xkCZ0Ej+vkT0PD6ET9URnYyIphNYQrv5TKuhtJxacxSqhnPMyhFeVxkSya
eQqSnsMn4/MjM+Njj5RPpuwKhT4A3yjX0fDLZ3Cj0yp19JNaiYeJXP6OADTDds0O
MVSaR7S5S8za3fClnGIsNdVT5ZZoEsWuk0H7GiA70VZYsesf5yJoFILQQ7lgRP4c
V48FmYFc1aClxP1zRH2mBhyGCvi7xwIhSH71X5egm+G9xPAolyonwxSAK/+7KX7+
Afl2wDoP+vvHqoVmNCHmq160zp1F3U+cQgLld94deAqTVkzmgkhHDAOrLC4eIJxN
MUGM5NDWdOwAqWNSVXzj57mTLzgmP8J0ImGH5WLMepV4pMZZRcmOPbG/pGH/OHZC
Zf3nK2PHk4985lTpavWw8yL8dsRO2qKHALy7CKZh2s1SXyQPwOTRsnTikPSwbdfp
LZBJqQ2J43axNj6RQeRauvDh8dUk38KZLRYL74P/BwrgMJk5BuFUwSKJp/r2VRFY
p/wn7wa1OpXaRWy7P0kmU1JELylGTycZvJBWeD35vUETTAJl9UXHzOdDlJQALiyT
eYXlr23oW7IgkRXVzwkr0vhbIiZpVhRrtDvzgQBdgNXq5upXiz9MzVPf/tXL/lGw
jROC7pRZF1ljyAYAmHpPd3Hole3Mhtwh3TRl11QmeXM262bdy1DE8ronAF3C0gBY
7KBesg3q/Swwg/tF1wqhTF62SCG3gITC1xx87wVze36rx3kI+040GNw/WKZXROSI
gumASJndkGC0nPMJ1Fzw1/MLQX2Rnb8zsnKKfSBn9Dffg3Kn6Jk4M8ybCmjKuYB8
0jSu3wIAH44RAM3YL3Gzk9UEx2oBCCrWJsy52PR5uVxst6w9bePWDbOS/W3bSdmR
T7XzFs94G7+QOSIxGpLaRrY3U62oxm1+rKVyk2JSpjTPxcsWaSvlEbjzyfh+C3ZP
zEcmpBq+77WZq1wFi08wfv/Smkh1Rh3NbCCi+orGlfCfGzNwWqMKWG+YjHWRR2/U
MNl98/oJbPdknSQ6Zcrz/zKC/Zo6bMtNPgugKwMjhKB6zXyphqo6FHLFM8sCO6h0
UbFm/ZpaSjYBbM094Ls2m3CVs+XVoQ1cG4iC4R8OpF4m9RZYSnrC3vYdK3xCld2J
DW1cxsSQ+sX17eVldA6wCvdk++/Arrt4uIvlA9OyCM/08tXSEHnAYr/9cYtfVG1x
NcXYpKQoWu1mMCNtLISbHjc0sq/LnfEH6fdMCJdvVRvzrc4bPr2oG5gEkXWb8Faa
odYwgFg6BNoto1DphCZ00EKixk6zG2oLooCeMRdaQbHsJoUKboAw0CJ14oY3l5ab
itX4Xy760yQnM+s0AeCp2CfTgMLz+gI5/CSOMrgXM2TQ/rn1xPEc7F/RkeoFTwZ+
Y2wIibU19sSEh+A4W43mxBoz8BEdPokIVhbjAf5x7sy0peJ3+rohHxGpFf8RHG1G
A6XpKJF6iQUhd3fHBqIraIREkIV6c2lW8e8yevaQ0JLQPv6+D6xhVC3C06d2dOLv
5MURfWKbUcK5ByXru8bgoxi+96q8CZyc4bHnzhSLZH+C9TqozlARhvlewhBB0u5h
CEjeg8lQNQ5c7f7C1WdNxqq7EpbeYRhYN6Vzo/FzG5mzzkhRnD6emRViEVB/KIw+
wQaQG0HoyE7EqahuEtOQarOedHpFhr947qJEbJFgyDGCrcZtQGnLDDqqmnKhn60M
O/ygF7UZQ9ur1fSsEQcGzEMc8j0UU/vaDAxlxKzSkKoxH7X1cPMeW7QgDpb4X1cs
UlrCG88LvQaAEDOQ6l9+CmwwIxi67tazzeKqL182D5LyT8Q5FqRPQ1JD9EELHrGL
StX9kt9MQRxEs/HAMKuAqIr9ndPYGgXy6VJgDZSebOigGLlt8U+xCGPcfMyvg+D+
pMz0zjTNSFF+Am/65M11OUiH55cg+XB+YZLTciRKNEoTZnVBbr58fa7KLag7C2ko
XmMYrs36bBUwc78N9wFsOaOrqUaWk+VTenol2CFzTrvOkYidNbUHgj0w3R+LBowO
96W8o9v3d0KO91UV/uRU9GPRGCVTa4O5f4MANZ6NNA+QrWynISZoBdfQYGtuL6cc
GWEKTOGdTnaOR1roBzCuNR0x1d64lUVq7jzezn0effne2/dnnjK9Biw02RLMClYX
/pHTDIm3hBNwA/6btL1MwiZvNWA6Abp6PvLTtb2kY/4cMQVzSwL+hXqCPp287bcu
mxppy/dPMDXW2dbwAQNjVDuqH4IU8kVqY//H4xX0sXnvluitm/tq6e+LsMzcgyNk
cb2O78lm6UWAglQHz/1ykfD+CDVDI32gz97uDdiTN1shAaR85V9/XQQLyzklgLzX
TRxie7loCRYKboC3YfSQfIZIjNiUg2tLNpRO+/Urq4dg1PLVZnOvanqfTdoZoIZP
+V0ztwx9JfD6jOhvhFbBVq8cK1OSfCaszkMf/OpdQ/iY82a/RxauuSMzdYRUfTuN
wkKRaHDPcSY/UcPQgxnvUPK+m92jEm8nWe4XPa5Nnsab0PztZKgQFBryaSwSP+aS
fGcItrT/LKHfxBQz5qHvZRysaJZWClSwYdFE7eWsoNN9wO34Ga7CBJOyOVtWSznr
7UeXlS+A9h4zxa5eF0D8omwzhVieg0lx0vuezrXw7l1dIG9i4NqBpVuhgwkSBD+5
rkXrwBDEyW28tR1olT46Zf91iRkTOjcX9PzPFy7LBwAx+YRX/KarpBjqqntG3eIr
H0iw+JFlbOnDc331ybpAMn4Jdbevrxg9pCzjBN+BOjk04F5swr0nT+icRNsEvE94
a6rwjD4P0Pan77sfcGlsrriheIW6Ws/EdOrO5PXHvKrgC6L3ylwyaJmSN+kF3qNu
B+3WjrKvrqFaoBmLzKMxI4nPcL2pv2gsOsjVDuDdGHka1IQ9jY734uFz2JKQqzJW
dNmGOvI4ILOTO81AFX0e4xjR1fkuoEAemTkfWOBq5IyCZssdokHfKQHirvmo5+v2
bsxezmo+IY4jIfyHG7hIsk6DXlxWCe5ITZM/pPsjzknPO7UpUAeTou5DaJAGKTvl
yESZABsjOU+F+csHfS+78xplExwsDZdqUlySFF9OUjTAp+7PbhvmMOtFoeSiVaGa
RdY1fBpPRLZ0qQUbun5LAJFZQQXG3opNz1rACSPeNTXjelJvZ4ymk0wyWuS3DiVn
UaiceAKMwOwFYPSme+tWj14N5rVSY4hrUPProCAljbi9Xn3dur64uJ7etU4YX0oy
8QsbprqN9kea1XFX9a60sc/XIFp9OXSB1bBPfJfTcyCU4zgEKUt3PDLmMPkl5z9T
6wWXTgR8VYBwPGx+WUlL0NA49/Uz7Jey2kZCInJjS7tdYBZR9cYpTxsaNrUhDGCk
gf2qmPy4YhWJFf268s8/Td5+Yy+R6it9ozjD2FFcf3wfIJsgFTeodoG2SP13XwyW
vcETWfPswN5fakls7Qh5Uqgwcu+0poBJEoY4DVoX9zIZvvZnrC1G6QKopOgymr61
Ug5sGDTy/PXGmdc0EBaXnunVZef0rewua1JShFsU5B2JofG7I+bWcQZntt/Jf5D/
/q6kKbFJY2HNbRsVVorp2QTni9dyT01uEHlcoAXoXiGtFRIiqdJFZSVQaXahTQ4v
PoQnJ6WEABPAMzLRSlrJfZ7CITXRa+6Q536Cqtrguh8fED6QVbXZbxm4SAHz4xAH
JngGEvaGh0TzeoqJleo2u/kfuV/ng2/RpZ2kNkcbuS5bA60fGNtb85TZqKEeWfYj
5ixgg8ppUMWm3lEbaW+XRN2GvcsvLLxEznHgcxfLi0c9MToTjLBGdkV+lO6iijxz
mCxgni8TouFtwJlHFM3PrJjQnk488ge+7PuSMNqAMp04x1JZ82sHHIHqe7engoK9
aMWPhqDqs7OQpCWkLlyX9N3kfgMRHg0iGLnaSZHGfIsuO+cvw4JTFw7kzGruPE+o
+StAVpiL7uYgNhVsxlOlNVy7JUZsAu0kEkkOS96LnLJdmRulqweev8Od6lebwjdb
HoUMxKsnhaGtCm0EhCtGg36dJw19GziiVxlPkVZBEb3U7nT3EAi6RL8qu+wjpO/B
upiXe7O1Ahh+i39lOLbbOi33W/dVBK8M1ZW3YI7iSI5UyfXINPdYYTtqtkoHxmVK
tctXka6+qk9ntZadirPxdOglh5ppdu5Pj62JqmmZHE4j0AFcNlLj5HTTzyd1S/It
HYGikd4/inalvEhWl63kRTQEdXiiwI3CmjTQ/Op5LZuK7RylYw9GRiuBWj7QTqDs
2X6HenOxWk0AsxjE0Kv+OoHXaII0N758++cCLJAbLgvwvyOWG7NJRAtWOYJbEsOj
G+cw6nwbjqDvy+X7lr4UgdmXl6pIuKnoMbtfrOtDfIc0wP77wyqoiSBHNqlSSs3P
+2lDIlmZVJdv93a4A0GtQvhLSz8sUQFZB3MwmFqarFum5wJgAvqvBoFXBOvGjybu
qw7qh1iQDOeb7YQ8kSxFVCdwjr24u484O3vhLq5QlSDgt6CtPs7FUVSj8nQjAYo3
kvD7tjKNA633QuxzLOXnycJBYZSwiSK+EzQERFA5V9GM07igLZF9IQtxf0JVbYYc
P5qwUMCeIIXqVe17sXkyi9reJGxS6GZhDTYKp0CDiEE26t/OrHbrIQWXdF77ZVrw
FSKAm+G1W9NZqWI2GXpWZTpQ9QQcIvqZgOuhQQmw7L+ZAfdA+5t7kD3Y+C3lWH6X
QJ1jCR+R7+e26KFKD51PyBZr+bcW4zLi8CZPnKUs0U19Y4RCwgK06JRqwLQ0oZfw
qkSBoEyPa+6Q6kmrYM8chFJu+iDRjCyAcqWK9o1DJIt5Whrq9G+Cxk/Rqs+ZtcRE
xok2mok4HMs0MWGvrGWiJYb+8UZcPGM/LpysrNQ9aecU/8hv775IE+j+tZcK1XIs
UElsYsw0CxT+nCyIa2tonu+1sw4nlsYjwsaLdW9FJ0obU0bEA6gmSDrvmk4awrq5
+NQcttBJwoxUUW52TdmRs7n4OkcktNAIBUFlvVyLfR9B4ry0AT2CvUF/cWUv+G/3
eVrUTh7hkPs6u5ZqLD+JB85bF9jf8pX4xrysiV1oKjJif/YcmMTdrAuRbaOnhexA
jiVk7OAaUhpyxG9t7+SdAc1rkZBZzguT+/nsdx5prGNj2Aqbgty6A/5vRoshfd41
xFZHhk80O8G6eWsn7eSHI8rqcJuvNtsGaeOWZNewB8T0rA2i87qeP2frhtGSbTzK
BueoX0+T+545f3OcnhNHQtlSOkLRjXBMX+D80j3cVgAS5LhxPds4QkOnt6qiLl3F
vp2UytQGv/haJhd+pdgW4rR5MmgA3bMJsDC0t/gcFJtf4foX40tlTK4pYT4uNnN2
UPCKVXcDp/jumNMUx5spTi7d22+F/lNJZgaWUVTnrJWYmsuSWZX1DNKjpMRd+aMu
xC7RjsWw64RxKyJodVgW8Bu7e5ktyl2BGKwom6cfIV0SQ5FdN3tVPjrUTlVKELD1
nIKOOP+O7ZHg0H2HYZVESg02YUUxGXA+b4NiT4orlqVEM4n2wCPsPvuDga46nKmp
r2y1e84RKje7nmPU7kSZpWNAU9V2MoNAgWO0ZGUgYo/0YYwoE6RnOd5uqF+Jq8+2
GoxjX+N4GJ8aB2YVw+loYiYZ2Vrt5XJPsQ45C83fW8MnrjbQFnHPFpw0bqoHF3zl
jyX0ql9tEbkCNmYjS02t47G7pIhX1nR2SGvKDKQJuOcIXl8InTydejH9oNP8vu/M
RckWwDXQJPnGZdI/ZIIY3l2z1U1u8lgPwHEriCaGaDHMRDBwQ+6jfj4iVr2p4ZOs
zTuaDGmh7Dn8CID5ybgIHsECTElKRvuB2BpR8nXg8MMHFwS2WXzkM7sPh9U1R5tT
bkuqLxNucmswZyp4npcbTQE67CcHaPd3S7icWGlFu6tUXudZ2p845PqDoBmglPuu
Mbro246ETF3pLmBPQT3smmgedC3i77pfKzHgOoooqZ4fo1GsNj2iIJepHFfnhEUE
U7y5F6ptlY4+QzpMh5z/T2nbzC28LVpB1uDxAL3imCFXtJtTkXugz8fge3vvtmhD
H1cHKbjYac1F558KL/qxQ1IBdGfRdgmt3oX14Qo7bmEICAyVo3rde3r+EKV8Di4q
XAUAvXb9qkxK+EMjKV06A5E/o6G2rzFPdjAmuzkTzqAFCEPdrojR1mz7VS5vZIEY
4lgbmf2hR7yLJjVgIuGei4/lEAjsgTWi4OSR1RrJHVgJeEFEGQZ1apkbWdwNZQxf
4e2fw9Lb0Ape4HYf6buC1cZgkbKoQqMjWB8NhnB+nh7Q82/ygdHTSqZBAeoIWSyG
ykV3yjWwv+gOaDbOd639fW6XImVFJxhQNVerCiF/Dm7Cg5C99EvZMu6QMfo1waxq
2Fr93Jrt3RzBYCFz0/ZXhfBo03+xTyKZNlbHT4UXDnmhd40jbh5KWsQhH93+OPCa
Oz4BDCAzWhRpJawjkvKF9w/iyzxEtwaqYZpewKx2HWDsCrdMbwzWh0kb5Qa+XLE2
wZxxqOqkVaTWZbykpLJjGyfSnpyasvEzFsSNhe/yfDl3DX0XWuWQmOr1f+W6R559
f6HUa0AIcnQNR97pEq9lqADKjgzY1plG3gkpdq9yqlJyKK0oqiQqOTquy8/nPQgb
Z5NCuBRp2WxuciNruHCa/vXBHemGQUSo6AR8UtvcY63JJD/Aa5rS62JjNDUoC+L4
U1+0EJ4+GOfxr8VTD7StEdAN1On73wTV6ogsl4BxMZpSXaLi/mwGe1wwNaSKphsB
5OvNbf7NTRUV+vdQp3ZTJFKj6wBzYkluhzLOXKGJWn+FF8kaQVscaK7EeAEbPQNm
OTcF5v0ptmVuN3SLOcBt1LNc9SGlYp+MzqrnZGvN4rlaX/yG0OYymVKw8NdVNxtF
inRvjvp1umwb4HJxPcXAu8eR47iCcJe51fltEo8oCT/5sA1g/gzUiNyhexi0nPdz
WMv3xz3uisCEjKI+E6A4z/Uk/sUsH3qiC8aWS3TCtcSWWbxUDzo9W5Z96bcunuby
X7HjV3vMreIP3sbMnqFzT61g1m4qI61FUXvqnLLLrTkJXs3fO+bHDHsBNdTk6fAR
GIsUzsgfUbkZL9fmax4Zdlu2k0SyTDJugMAuPy4ZmmFWvmBjlFiSLEo6SqQtu1FA
o73tebV6q3cgadEbI/AGm+Awd5xhSKEziBsy/zIsD73lzIx8tuoZmkQVrb/n+WuO
LJOku2I09S23Zeqbe43Mfu6hAnQ1iY6Qytq/6HPm6EsWalOH1uruwy6a1BCPcV0x
JxpY7yMwzLelWfKxlYbIN2gqHJLdAY9nwXfdYkSEnIEvXKHfmn3AryMK/L08FRwO
2UI4eWOVcUH2mKU2SoiodkCAkwzSNkus9SYltxjjGY6fSAvKjeiw6edtH14YeV+u
IKDzfLuIol1FpPx2jVxj+wdgqsrSXyhZcTG/+SfgycPp/aWNINM/krtGwroFdEf+
i+3SYoRTGpKm5MElNgU+RSizLrsADuOVi7K6fwhgnAhp5NvlOfyI/7y+taKLjSox
/EmxybHlIwA8s8c8ahdBksrr8lcSrPipW1puQYYoqAHXMgYhKrnVk5nWQPuE2hGA
XNFG8o4Z3Lq4Xv+DKWYq2w18VfL0ekmgeCfbhoEMsLeMlPPoNiDCCcg8Z9AXcYgC
vjr8fQvHTr3okEk6/4C8zwDEKDdCAyJ1lW+c/DdczHa4gqohmAKaLs3LS1DyFZl8
gCNRfO4m+f1TadHi3UOXFCiK8DmXv867s1kRnDocv4y8O5d+fimJyK/SzOExS+s2
o4By54+c4Pqab9RqPneys9S+op/BxjemI5EfRURjVn86gYcjGPW2EbK4KzGfZmpP
92OHtXFR1SeTK7cpv6JAsmo3DgmTZps/nczVp2lD4trapKgK7zR2/kb147Q3QEyE
NwA3zbqVRBX/nX5jm94qsanb8Jzco9vJrfAP5JPOkI44dnNSH/ooChttBH5RDx8S
ermf6uXoYjCPSPz4TPErGBNzqg1A3+35HonZUK+sqfMTkUc6sy6DyPfyGvXvpYLS
9bydquFsic//G1qgYrunn6wTSFSIaXOOX7BcY5aH5TxuJn/pd5C0BpCYR3dKqHV+
hktaxnuQMZpIjECXR/JN569h1sLFep8q3nV+1MTl4X5Vg9YZP4sbnn/X7F/Xuroo
tcK6jrhORrw2m9V3tCl35o0d2pHCH1akXZuAoh5L2RptRtgqZp+L9KVP5yw5ZBYf
NoUMlrEvHarttOA3+rGrDCA88z5b8kwy4JpV4+DbyOvYHssjz5eJ4+FBvAiz3wnX
4pTXPC4ZoktpgiRMEmwHWSSRCcJ28S3zz8FIS/QoE+qZGBNp4BNF5+qD/C9jt514
Diqjmp48FQp0LJWu2pT3nClnD+vGIvm4D+95njm7FUdns2PQTr/aE/C12OflAEaA
BpGuvgOyj8ZUv0SQei2t/Ghlryf4qOhgfIn9PR+SoEWj1Oo58zfOFynXREQYS19Q
1G10t2jjKXYNczVTL4VxXGLxt/dtRgQIyv+O0vdfPgmHCA6u/LoYH2qs/PYVKC2S
3DsWQTqeHYZUEkfKv4BdSXn4wISyaRojNFpp1WlD1fMCk6OHJcrd63lJ0Wdkd7KI
nQN3IYt7/aB++MuW8xwXAn9KfLR5dl+K6zjsJd+5xkCkC5A8MwoneLsEl107nQct
qovowfyzaJqnXhLFA7TJ9kjsR80jOURKwcvlzMxuxWyKwjQdIZ/ZEnY8be4pQHux
e+OKg5QpFAOeBqiAXQOgPNC1M/cV4iQ2kUbyJwscPTQRdmSdTqyoaPi6WKdCQF/E
QDD7jV0ZkoWcPf+kWOEKTQYXG2YAR+R1e/B2r373oLAHxzI/+vilRFskxu6CCSVt
BxMqSIc4RLiC+BDcF9f3Yw5A0O+vnh1pbvExtrScrd1H9cYW99Xf3odentQ+P8U1
BC4HiZazw30fhT2YN1ktb088CNHdVzrUF31R/EHBrKMnztYCRtssYXe7VRmk5vFr
XpI8107+5lsXdbe1fMHkJyw2SP1s9B/vVKU/oQylKldB0rM9enMCNQMXvaDnykdP
D6CddvUy228E4PSf4ChZsj13giWhhBpspBFIdEQCal0fBDrLzWGekj0j07yFBX7v
bG741LcXPApVu6hs3a0enilYskg66Dhb/yn+mKcMl8Z4kg9waj/yAjuGw+4WzYkX
ArFiCq0GjNx3u31Wzn0RIWT0cL89XnXpQ6uGHpct/YHZt1YJbREEqxPAhB0fR0r1
vyAdBBy0hI7i5npwygTRo62A4+NpLhBC3Xo4kG3hp2mlKRY1lkss20Otb7xOAoWd
Mc/F4Y82bnyqDar3dGNpfs8hq2QFE9BeuXemKhXfjJRQ06DFZTJCvKR6KzEjA2fx
JZiKuZFKH/fhgQYOuW+9bDBDkjvmDEx1czNs+oEpgTM1S07BYanbeDu6ktfYvplN
BMN9RLcXHy2Ikz1X9I+f5IlqB0N5rU2Yh+Ig74s0aBbXJ5yafZdeW7S8UoHcaXQb
cETp6sOAvxfNub4biSJE4RJ136/uNeDwAxmEIlLsR38E4niIxQY1G771Vl+q+/8p
AAqj6I7BKZD3UTD6Iwq4qGInDCrH2You6NgO2al0pkrvCFY7MX2EFzj+qAwQdLpq
hyy1X2jQsWect+N1CQvEcVUEG4t26nucUZ1Kcv5v7l+fNa161mWxwbdCGeKoVWa2
a+TLCcXSmT8NPh0jAaAQzPs13Ddx+DVXg56nkxYXilCwUIXEKx4dZXuY2hLwQLjd
l1StLx8Eo/MW385IvncpSn90Zc9jbcwvZtl4bG2D6dIuGOZhapSHrVQYf2HIxZG5
RDO4XvqQZvuvrlPcEKSlSkqYQRLa6JZ1UK0e9MM8JkghIcfXuJ6ThL7U3mMfnci0
qXuW80O6nK7Rw2GHUW/FqlvztY805OD8j1gA4o0i9aHEXvfeDLhPu7tNSwVkFy4v
X2cH22phWrgoVKZx/6A1nC3FKtiaqNqmutMJ9oITRk5YzLd6I0mbHdq+SYQBPRG3
rKU/AyOEfWe7KHVg6eZxYmBStW0pzdaqFwC5aZkWDfY8Ruc3LhfCEr/q2AnZOTEA
rQ4FYBboQ5l93lBgnoKOHkjsniTGvrwRMrXLOEA5LmZp4ImgRJs89n9+8+isi9ok
UAKooJuAXCy+MRs2NK2zTN7a9H2Xn6vWcYE3pBihhUkTSVmIZUsr88m8rXqkF8Gj
cq0JXhth231q1BzyQtFTlO2qOtnRpWiURbk/IJxmGcRfVhyXnfymyF6nKdLWd/st
Qoy5pY58gSlNV0j06s56jodFDjevfTfI8qzZpN5PCIYmFHIg9bwPeJ52KG8lmyCH
27zIVwbjSd2ZTG2Dd+67gFUYB/AGeOf0zgXCPUV4RtAP1FxLFlDi7Zo5V1gc8HMk
p/ce4vx13K4GDiXGm+2sjtossq5XGajEJHATcZ3KFAWM/0NuF/usvielhhv8y0b+
2SMmoqODTPs1RVAl05YyvOPkZqJAElxg6MX3SsGq6y53LiFH0UUIwbq67ZnEgqGy
Q7qdOhh4EkeQlJnJHVh5VUAAzlZU42GsIEWg7BBPlyLmm5ANl26rOQ/wOPsJkyPg
O2BsmncK+eoR0TcVTnjPMq6hZm+yppYYKyF7IB1m1nx+Zk6TuMtSC4Kly1DyNzJQ
LiRyJuLmj0IW01rvFq163h1AsZSw4T0cAV5NAdWFE8j/szH7vE/FwQ39NzXi9/Sn
6dOs7+yjI4rQKpJJ/Q1pH89kbjDFSzSF1M8eiTpSWe7KozRQxADg3pHjNGm/NKfR
FGH0kMw9MCcCWbgC2G3FinHZNu3zSMNk7hUHeG4ibvzwni6P72SoYd3tGS4Me/uM
KOHm/5OUtzOo7znJq29c2IwVwMWixrB/3e4a7H7bzyuRpCOQWHU054uLKgZIDE+o
BlFOnXaHP1rO6BnuVZj74fbCABdAntKt+xqC7In3pTPXxYTKPH+T3pTm2LNJWjfU
oRVh/++hIsxrov/tYHf+QJeGXCihp0b+YtWZM8egY4zRkaFLDzSmIKqPudQj70MX
UDXEwRELWffsMZG+nuAwgrQOh0hJcF6HdEw26w+ZYkQCVLcnkxHFgfwKQfhG8OSI
mhR8nA1++psPP4SKK5Yfa4V2odSg8KN7kOYJwO7j/mGFLcQ5s+sCvy25sh4m/BNt
g6s0XcVeCXgCazmn+FXXwV57BL+MBIeAg7nuOEWZpRwYSPUZKi9pdPOwiYyxYHyb
Q0HBZxNBPtpFTpC7DAQA+2aXfP4HdGKU0ki9w/t0zxMPeMLirdGKAwnZbi3Yin2a
UfrdbFqoweg5oJalS2aqyCSzcLfle6kZVzgH40ERmKURQxrBw/60XzpbljFb91PG
iqMk9uS/ShkAPPjFnpK+vkHSqX+WYKVeMNjmXox3cEla+869EIvTpy9auU1kNaHe
wf2NI5N7a/QCHdjohVOTtZUfhAWQ1sG7+qC+KYjdRgCAtAarYyR7/+CtjMxp8dYX
CvsV4ifJoe7rbCchH84+Y/s7tL29ITgy3ris26GsOdA6OVvAyr4Z9ibuD86rVhmP
jckgQBrFA1nhZktVYZVvgf8G+0W9YRd+l2hDosP+Sq/PZwSb8vN05Or0GwLHSOzL
ZLewIleMuK187vayKK/mOjgzkVSEOoeHucUKz4Q7mWSrrNtRIfCmn5+I5HqZDYxg
kkUaHjiXHlnMA0/FcOdQskLiJI5f+NMTedKU+dimBmtQPy63iTPjMfvvlt4IIUq0
1oiv4EiuwF70bHOsNnXNaTD1Yf0Az3U1tcsAYqDIdkpB2OFhdFeNBCKl0vF3mOiz
kY9AUNX34ZYpBjXUlM1swlngOItDXadXvdFckRChYsFH8XV1bo0WUdtKx06Py4if
Q+fm9gQkSl5foshVMxFhYKS+ygfHUfmPF3kPsGo+/ICLpw1ACkt2O5vEDo+HGMfq
llmKhHwYQpD9GsbZ9lgoJgYwZjLVJchOQyZdcAfsKQhSooyNdnoUHMBzIwfrwKKh
BJ3/Op2gMNx+7LO3mjOUjOSvJLQi746dx1WUfRpX4suGD6TiKUYfcHLsII/La9xo
/msSuT4csq9sRqvuAnK0sIbiaX0DSesBSUgxsUZz0PuYSu+E34ExbXrQvC9Xf2Wz
+mfR13Mi9tjpXKPkRZUSajDz0gPdTuG4RCnxyDyQRgdw8jXF9YPTaFKduWUok1Bs
lUkX1ImxGf2C+T/TElHkmPiuA7r+wz1nYJOa/Ha25A/SSJgG7gKEg7wGFPkGr0AT
IZGMLXu1eV+i4YT16MekVXwqXiu76vbxRxYZNHfRcNCj4dcxiE55iLIdrVGQl6oQ
xRKWJWfI+E7uRaYopxRV/6499HFaqpA6TBjbqNy1PwMRINp6+y87pNFfQV3J3YZ1
rDQMMhxzmn4VsBZt1lDyBE6J/Fr8/e/BaXgvuHRLGlCy3Nthv92O312+Po3EK6/2
n9jEDXKuMudieW/E7w53YaLBut3wnii/zcv19VPICJ9h5ofOWsxgcW4kcvQzniq7
xcuMI1Yev/oiajKkhp83UoLdg86+xu7uatRJuu4FeBVgI+jSmLUessEekA3BCUFa
HnzrwqRto46+q1GfhJfAfxWM6l7opqnZ7lBERqLXun5Wn1UG3CfWy1Tn5AoGCyRF
LTYt06jlGf2QLNTFBsI+aJtnRmAIlnEJABv/TI/x6mNMPSj0dbppgpdYDsKgsyQl
RP1F2DTj4rODe451UI6NK6slc0Fjg1G+41B2xKAazrNLkHGjq14ds9WYsx1Ukgrg
gU+W3vRP1elLD6mc+P4GIIICyElOjtGtZnskHdDO7GvcBCcUZ2LfqRIbypMpvL5E
3Zt5ZSUyZhMWWx7rKWc5eYUh2EUNZqaXZ4ZZ1XeJSc0MhqRriGiwz8UCCrDH1RfY
nqGCqAPy9YPm4iiseoWNzH1Up1ankMvHHsLCI7f2NBRe5Q2+XO7umTTjQNh3yFqU
JNxWXNsPEdD/MSyFwK47yd6R+9NFPF6B869tGWNzDkHjd0ScL622aNDzWaBExN0D
r6rfFJiMaN7yBy2xsnx1Un7AMCX32WxIuQNZqHK1o4zEEi5CNJhotQ7si389mc1P
y5oL+M8m2rc1YU3pYJlCOcYDZGb7Ea8O7EevWPAe0Lp7G9hJ9ziGjy8K4+vQeIYl
83+EQe890mKwgS4HJ+jGzMcXQ5OUgxKyrvxR2dvEa9Aiki3ugTCQkgdQrx8NN0vO
rsOmWSy18U2vfJFEfRWZQx/LwjA2AFvRFYt3N6ka5wIqDip4nuMfWRImZOx0KMwI
jy0vsDFRAKrlOfJdPtSUlVt1HwYUp0fwWuKHl/Ts8rQ0Q0NK412Cb8y3Q+qoONOY
uZc+Nlq4B5O4WK4dLFK56gz8TNUiXj4n/cSQZWbVU5Lm8uGBxqSRO+JctI9wYA3x
CcAxasH9IOypHQdmHiqC3STMXFvGmfaPa/ksvAyDr55Wl1D3XpCLgAw4OqFecsRm
irM78Tm1i5FYjYWVKCi2oI9dX6xLoId8QVB3XpdLdJuMwWsHxLZcYx8QbUogSHMY
PyVD0L8TPZ+LnDQ7Hfsm8TgLy3pXgqz84ZSpPfeBCm+2fKs/KlYOYCYLi6cwkP9Q
beO5j1G2Ts6vJOx9Q7qG+RLXitvIwKqwG9WFFbn1LF4RQb/UMp4p796niyanOAbb
9eb4cih82sWTjb/n7NtR0ayemrAMRJ/6nTG+fKij5XX9YSC/beC10qjH6Hdw8a0r
on9v8VtNwPDEMNY1YpU4HtW1tGUJj82A0LLzNUbaKiOcP0qB+vqWDe8E8yBO2swR
sCp6olGQ/b2kAntkdNY4Ry9DwEsT5/watsBM4fw84ZhchETXkHlhodkv/9TDBXYm
CEQec9/6KzHx1mIAH4XUJYMSQaNywY/nUrH1lTFVXG9Y6+OP/eNZwmbm2LwrTAVL
hQ6vHIuXgAkwBSGw1kAdW3dao73x0AVV5xlpGYr8lhLm94iT1VEw/FbvScxyAqxJ
5xbOYNeOiX4X9LLFqlZz49fYSfXlx2XEYKrIwMDZwgzH8P9szMfvQ43BMs1NwZBY
Zh3cCd2jXH2VndbrCIouW+pdWA7i4vJxSFu8jqr/g/sLRa+qD8DtvVQP8GS8r5OF
NQLEek0/1iFF+MBXzPndkj6dwusKVbU9QS3+6oljcSxnQElKyRbHrB9HUgJr9f7v
GKBtUn2jEAl7Ah2K/y74isjgq5ifNoFD0KogV9jlzlhl4FYoscInqoxeg8oHAVYg
OMVBuHvp/Tbyv4BKo+zqxsF7q1XZHnfw9s34sc3PDH2jSKj7yLAXOlrk2LCLV56J
T91w6d5m4hjFfTlQDQlYZzX7ixoYHPG1LOUgm6bYfNX25ONOnzNObIfXseO7Yuhj
pfRefOOgmdZynHaJiN75a80m68K5nnvshYYsc8DplnXLiPDxvypnFVNCAQUD6eDn
6KQd13GpMceQhRdKfKNbSWN25PdivdbX7mipNu7eRHT/kvtqvRbWkr8lF+3ZnCeP
Ia3p4d9NDSZLd5K5tilKPpIUO6FwE31yJI+CveJA5SeqNkOzTJyb55y4GXfcQ5nJ
MXfYHIVemdGj+tR5Fdd4Xasfa/PHXxpLUzXOILTRUH/fJaCDRBVdyUQxRGobs6Qb
aM6ioyWURfTm1f6C1yTl25nnHI+DyX43nstUsAAGrruM19uyLH5zDP8v/CM0OXl9
mlxXwulMjZNmMPe/VONMlnAfqPK1Y3YKG8qyC2XqAIwetiPQYYbyuTgTxssw/Vc2
F9df33+yP1P4QVTHs14yYMITECS/KJAal2E2X807JBCLe0jgOfopL+yhUfH3BJ0w
v10p007L0wDOhgkZoXJOg0QOS0mYkZyz93HmxYl3QZJjxXAOFwJIno/wouaJE30T
DvkbPfNoctcWnUCROM8AaLogzbQKSSqAOVfWjI4wgiAfJxZg9HuntagK3YuJAKYj
liEryfKOUdj1HIKvO54QR2Ti2pvPOK6GSc/WlXI865OLXwMECeDWalda4sbmbOFs
9ouqpBmmRGllHT44DOs1x7t1W4XhAgi/vjMS9Dlu6yY/2bo/J/vZQNhBUu/jSnqx
LkTsP6HV/THPjrfRoTHPBVN16IySKpVDoGWql3G0b1bLR9eUM3qB1h28TXkwRWlL
MTh8yz0A2dk9dhOCdelhp3HZwizYpLKiAS210dTevcIVQdqaXOVEj1KYi7XM1QPS
ykm8lpnvOHxeBtwbmDPgH+tmMrmmgy9A0kZYKCtk2M1MkWzP5syHXZnWf8VquL0c
S2JeRh0YtNpnr2hSY22ZG5/eDWXoTBbXUEJY+oizyiG8pNsc/EphPq+aiFYPZi1O
lLcRB2dt9fR9x+xGDVwzFCgE325Y0q2CFaiV7pGjm+X4QY5cOoymPZrtBrbACepT
ENtoJNdhRIoYZkINuZgZYlA/AK3yVRjoNFANjj8C3tZDdZsT+mj0T/bEY1whcwxB
3O43nyDheHVWU5lzIKQvXNLL2//T8d1DOlPKaB7HB1yAVHJY7gKYIXZIwfIha+rp
UawRNpIG/SF63meHAydsVkBWchVNOfTJmfq+lFDHenbmIEWNzszII4E2bNRQU+X5
W6iP+n3NzKudtqu3pl8LGk00mf7uiY0Vto2+Ebn2hW1EVycyNqCd3k2DDRtDsIfZ
q2vhQJTPOcjmYJyJcJ6TiWh+dL/lOWd1Lf0EyCXugIKSS3gEF5vrnKuCd+J2imob
shSkOP5b5UjFhakJSitrHpZG5Ujlxl2c+1yiC+aSD1/Laol6Ms3Y2oUl9rxv6+Bc
2jHFh1fvxSQJ44rS/jMicPL6EZJ1wCBEm6xb78SsAgqnPt2JuRc+sz5x3NhhN5cd
E76qLTZ02ksAbpPqk3PDJdxgO0x94kOZOLgCK4OvGhscS2+xTE5MiRClFUlMvs05
o5o8zwym4nBTP9/V7dTpzlRZNS6M9eQPLirCilDgIW6Enp5CfB8dLoA+yDs28+8I
0K3nTZY8FaEM3AF7M08EYIK0ui2KdsvrbCu2rBx0TpGXha07ySgZ9yxmR3VMSyL6
DibaMznMdXyag1nSnJxvAuASbOrYReJg3crq9jxVGpNmG0waRzj8orf3wK5v0rKG
VZSOsdqYq0NKzLK+KI42v7j9Qx+EcfacJ3Q0xm/HHE1UNrVbbNp5nP8JDbXRZA5k
bvZhtUVffMH3AoISMwzUyxw4hzjTfgNdP/teXyaqrqCS5hw1EkhMpSMWMc7r6KeO
fWVlOV13nWFSQ+byO+1ebQy7wf3TdleSAzy2NovJ19wJrK84tF/jHHj8v0VPkLMF
zzkjIYIlXWWPIqwXGZSrWpplCKVXeYGFPdZX18cPmbdorTEhR7Cf6hXasXDiCls8
84yrbyaHzQ6NM0kp34gukA32ITLuOm4MsXEgoQMFIzTv3HeKg+h1bipY53D8gcoG
LQCtb08TVWJQ9LIZDeuE3GGNJvtRYfIKNwaqK4h3pDiqfK0eMxLDD3ly9OelV3PV
9ECVjTJc7OB5I8Ogp51p4wg+HmJV3D/HbQ5tAPmY0F1ndUsAxBMSEVTsfBaJTdCt
1nrhNtMXK5DqcBlmjeXX1CLuBs9yyBpD6VLsQMmmA//nI9K630X8D8EgbXwdCIDE
aAqJfvoGJtfpT5z3N7q+iIGx0xqW5egcxd7I7085z1yP0QjAkUaRu0mQF/8l/qBR
E5cKAvmkEQnNgZ4A2SO/p5VsmSbampgm6ym5LhimeYdBmjAdxHj7MiKbmoc1KY+I
/+7MPda2oUu7tLCK663ZgHS9DJ48Ij8lu4zUXf7sC31CFLVS4oZzNJ6O4nKsb89I
oUrFztfYrORVMXttPwMCQVqm6cfPmSvb78t4FiIb4adqr5mnCc7tNAgp7ufgc/y0
fRPGvpdtwMXXVtKhgf4FsOmmGbPlsZzhVvHssm+1K5MzuXspnwubPOUEAGjzzMrT
OZbFLfBIVeOawiNC7HZZlzMrHecEeYPvYL5ADF7SHnxWLyIHzE28gv9TTU8Xd4aJ
jy2vGbGees+aoILKsx8YF2fXTB3Y6hu+/YGH+sG4z9YsbcrCLh4iFHyNrjBZr0Ex
nikLI79RM3BK1CJtV+aYfe5XSbfcHrxSeEhfTIN6xQiszLccHBO0TBgXnSx/sQLG
EkM74nTTPengIA0CDv57bnPgVBYnktdu6X8iEMhbblx/6vmOJQ30HAHh6bzAd0Zy
xtEgn/y7STnBVzLNT0gg4FFbzTbopq6mmBN4ybUdBRuEfB97B4I5KPpLnPEbe8VH
JCbliknMA4btHOm7yZeJHWnHjDCdtgiybCc/GL5wZPnPkGjbEsSp61+wGLpf5Bxb
L3Se4bC5WTMgZonnO7wLlrmUbCb5neNcKkC4A2CXV8eS3BSg38BZN7xcy5pkXEE9
DZ1mKhU+KSMr8/JX60JeQQcDX/Az2j1xBThRed6LE08hq/cTyi6t+2IdIboF4jfr
BYB4uR8XTM+s5MihIxtdiJ6afVglc2Vd6axjsGjbThTHsstyZ4H29R7Vi2plwyiS
vhsPWIKXU95XCHDmoM8ExuGLVzTsZYmCdHLCEHz99//OtpU2XtBveAc6K3o3nImc
qdXMCT9F13XhpSVBgF4wChq0P/2AunNyBxu/xxXlGbNdFWpxdnhTmhPc1DM/l/yD
IzDFFknqH0XPnEIx+pGKsiPdCybEvrbB1smKCNnaH2IW7R8jIq/5WzeIavVBc246
cyh32D4am6WASeBGj/MxfZ43eEQttXhXlqN8O7BMMfmUFDiI7LMaTxA4cC0FR0c/
A/DHRm9HX6kBldyJHNY1LDe89c9jxetTd9GaeCi+NqlwWtUpLuHex0eDIdVtr0hS
mmU7w1ixNWuHbf18HncEz+0sgdU9w+Td7ca7eQj7T75bfBRuOmpbI81R82eqbZGP
BwY7ScYLv1ZiazWUGPDK5hqgpJZKjUfr92jFHgmg8qDSqUkuxrgWMDTZou96Chbm
x/GOgcrTGiJ+SEKd+JtgmbZP5gChBG7s117sYHYRUkN4er7p1ohJL1nVEuJ5ja7G
jpicXubV8/sByYlh4tE04pDfWkjnKdtAT4WLbae7MApdEU8wBIpprzxs8GnE5Tdt
oYYQ7jqBdMpDPZ5vTSD/+70h5fl/V8bA4HoI75nrXrkGfNYLQjtg15yiKpRyq2xZ
BRS8xc7rvqCQ6Mu5JMqb0U++4Wyped2dYzOeO91M7oHHkRlHPMovLEmD8AvWqquH
lvAbSwtSDe8Z9TQQkQiPD0MgL0aig8VejuGfkuePn0cFTprdXpH3NOJSqRz0d85v
nkJQpOhSkGlXSVymKUJP338bIrPWVC1pK/KUMQdqqa/hZYBOzvizVqbUt9n81Po4
bTZ+F/ZnBDsoSQwA/b1HbMZJCTL0PSE1pallIiYt+aZt36OOG3QY7bJJqCgZY2xV
q/4vvIR0BWwdTowETHoz8H2WE+FnJyobZUJfmjKMMCWEph8kAn1fxJYqFGq61xk/
cK+xQPdY0Rmd2PszUYKn8sxO6LsjlStkgtT51yxPoYq88jHtbWZlTcNPqqPpURxB
vw54tn9V8QbwMFCjPEoVcxfxUK4A5iC4Vgc0RIleTqCKS34iY2/TEPmiNaezrfk5
iPwy81PuXyb6ozD/KHLyI8Dw3aeHFzMOv11mX89Jpht3KzSuaF0eoLwoG5X+50XJ
3WXnaUw92BGIIz4pBGyNgCJ014iem+oVX6R3xVm4HDThviTqkvYuJjPnHT1j38PY
gkcgzubG6ppb3egvhW46QFO4qthDsGMH8MPTjEJQKvPVxz6GCv+NvdgLj8NBDeFQ
M2plu7QuIHC2V1N2qGshsQ3KT4L3iaT9WhBe+papWv1rf+B+zbmoy1gjBsL+cNcp
p0tJWSg0yLC7YLwPSnHgQa73CZpFKlm//P8o50ajS77sJ2Qf2DHZNnuuQo311jUV
A8GDyrk3jD1Ym0vXryZG2lMIAraD0yOaV+/5qencVJFwbCDK6BflEbFpNHSzDJjY
fdb6stgNkekAu/4yPrw9qeDUuDUk/gZhZTcOFYD2dVSN54KFnGl1MwedTOlafEKU
sMfQJS3G0dokxBcFvAjjWYNHUojfWgZaOYaF5M/cjdocTHiaEtTW7haYM8eOtKyZ
cs1kjgajR5g7VyNKpwW6YBpZkcJ6GZVscF6fXzUtVfDXOXDFMyFksiQGgkVSrq5J
PmBH/Xu+gVxbgPhYkPyhQ8cC4vsyHm/FAaLqIwXgNCu6im8w3RCtnAUkyVZsYEOH
1BpiDztIxXZrxwGKpbnOQ5/9P2iaoAKxsx5r/U2XpykzzSM1nWRjJ/NDvAmryJp0
rNR7B4YT0ZF0BDlTOSPgE/Iwu6xPMXb5+GU2OBxGm7o6jTT1wnNntqDKATkaf58O
cVR/j6GZ+WipFSdMnTLbUzopPG05+6/B+xgHeJEfg2d2gRVkPAyQdDkaBIgA/JGR
Uw7KAd7JglaZuJR/gocwsA7JJazKwrO6XcrR/Y8IgeRJFXTfrEsz0d5/rJhJWh5u
C/PMOC+Oxcp9nPxFrInO6F00VFQopeTiWetWpCwNPYUpWeu4Ivw2RJYj77bYmRLi
L+k34KdD0edsl8qV9u/20Ms/K5M06ylY8PTacIPz895rja53Cs2nhulBcOs22M6w
vL+U1aVZ5vp2noyuGeWOJm7rl1PMTIOga9L8dbrfN8KWP62zMTSuGPH6ibewRmUK
oNIObW408OqEPgCUWbBT4VNUYX3MWboNME/7SNkKvifFI0BQLYKSMrb0VH7Bh19J
lEGkhxzz1m0ER3suKbU6znbV7VJ+64qCOjC4w2Rt9jv2aQEmOHN20UZgufIBEUr7
VgH0VezgcbFUoV4hdZ6Ag9ZR2zlZPpM9hZ4UYAZI6RuG5ZL+BFMw+FGWuRzZb6AL
Njx83Wjck6KIf7dl2CqIu9iq+OfQ4xCBvK1GHkX8hcEjHzZ1XtW4ufWuxQ2y9HjF
0vihax9MK7vxwDi/1ojog0gf8FaCTkFFOUfRCb8x1NAncJ+8OXMrRtfvbOh96L9A
7qNv6jd6JlFXY+6C8T/bA2OmkY5viwcu8GdxQSzReNWW7YFTywrRsV5AXzSsfiNI
Dk+aMSgav7unVeTPGvKADiVD/NeAC1ggjkhGNkNTCpzeHyQiUsmeR9hjgSbLA58/
X0ZSgsx0Xx9xDaBRdvRjOtFOUNELtDriuBBLKy8tbOvQSRxVHzYZmuRyQbkq/1Il
pzSpHTx+eusjZ95408XicM9p7KRoCvAaOJaOLLcLQspstUijqgc6nZhBmZC3LFjG
A430+QsHUho0AHTodUoiNGlBDKfKTT7ZC/y6Rqd5PFxJspbO3JK4k134UEWFgyW2
IfB1jVOpAHhDDTue7wDlPTokFGyJG1bqP0JwAElJzOTY6V0XjOXglPp2CgtavilP
FxooTmBadSInPvx22b0LDIHKt+zbfSbb5rxRr6XRoVoSOoq37Esu0X4zbEFHFC07
FBNgNRpkdQ48pviLGwNH5r9mP5D6AWZ2TjIhrX83SIl341DnLCNU+vzczq4Nfb9v
qPq6FpzIL9BEajaVWVaHdn76kZpvt5ntSUeMQbhG5DCWOThN0wok3wQDcBn4kQNt
a9dyV5eUK80b8ear9eu2smv+O2SM9Qa1n2FBItQVjaPT56S8F55gLVSmx7h9iHn4
fS6dCvS9NCOcE/MHVdtbeCVa4+rnDWxPm6MaNOv2xJmrAfQV4Sm2CE63McVlOcvf
nVTcgXFDMyMuJJ0ATKDPP1eIUOIyI+UqdZwGs2zrMo3+f46uhUL/c2ii1Zq/g/Ao
L2aMJ0Hd8StUUOxpI64OhXTBNZB3vVgzyMlMgo7gFG6EpXxVSll7lXA0Yfe/qE8P
XVm6l/dQ+q2CBycEK4yMgG1k7LyvMT60wb1B2ZX+cWA0XSE73arqhgwSosjPBbPZ
WKxiLjiDfkw1iaecu9RvWXCgg3tXsJ0FaACBUS3EjicFRBHLPWCqq3VXnM3UhGNn
W6ouWJSiozOl0C/tTJQjYlfs2vXQka+XIiiDtnvpxtXntjNVEjIQdR6yebMuSA5I
LXsxcS1CP87I7qcvYh10ulDMBvVIByFTAhB/eKqyHq6B82inOi3A76xz+pQ+Vquc
eeetPMC2TRHuRPYUew32wYIxKh8BbLc4FhWJu3dxWlRqje2ZWMHYNh20TsBQxgK1
CQSMv4dpfPsHodL8WGQiQhEW8eTE3aWhsUs7uAFTRU+l9hj2HzEDENyoJzRipxnf
n4oW1kRJOh/nJFH6z3vqBE8HhB2LhreYwiA52+a6XNXmFGAe+kBIDwZsUdC5hQUS
Wf3zRmmQBPzHhA1G118bW3yHELizoLdOI9litnC+MiipZzpxNUzEpMJLoGDKMRiS
32Ew4ue8BjOP1mx58eSGfRhyCm8xZ6zUJe4/2evIvcxGSJgSeV+g2l57BWLT2UO+
1lIVTbg6pLeVDQpdunEZiGmuSRkJ+ElK2yGR9TUltKXZaWHPq5vszp3PIdVHAigi
WIImZJViDgarl3imi9nBh1LWj/eRU8wmfk6n9HLuAsySpiszHQJ0s7nfwrT4qQ1d
0ElcqYSssVK7XBym6pnwtG2IbE42rttStxl7WtjSaZV3uI0JM/jxRwaCmGgIlHKJ
TgRG7/X6vvmLK0462NfqXYqftOOJX4o5wFduZqet4qRZpgqMsrprYX3ZF1mbGc11
c1cSCi5aSB5pL9S1OvlHxUDXqzUibtCylXIVVJk7R65ZGxlM9EN6uZeJGeyhwQks
A5Jp4ZONA7KQkf6UN0efWEA4lJ9qARfTl7qiRe9x65kamlzYMeHjn1wjJX5PIw/Q
UmpVRUiKL0LBKgn2LNnIVqnCHvkSL67mzRcyKu/i1mxLfnMnqm9Dxk8jpl5Ikcpd
LFDrOST+lr210GeHVu5n7iPWgvPiX3dRLN+0BXIDhB3TOiqW9ZFFH3ncjCRuMXpm
vLzvzfPvTbgS2I8LhHWedobNIVAIFjmKGsxuzSqhiL2XGmDazqcKy0Pv3YGl/Sf2
2QoZQC1i/pCGaLfbyuUNBo21GL3SUm01ycwdxpg48w0Vt2tSP18QRe9mUKgDlMoS
XJgoCjgJjMfZblSyRztsiNRKes5Ei3XX3wS4lR7icVX5oFePtf9dEsvsSecHUchT
j9lz2M20sasxKMSiIHZEdjZGTPN9lVif4Qd/Ty87Pe9nnNEErku0ULCD2SCRpn3m
a5/vub7FfnLWrA2MidZB91t6mZUSPGIAriHIz3Iscu4XE3dg3WVj6RxOtvWpR0Iy
Kyfdipf9U85RkgxysjQok6upP/GFvPeBJ5NC0BcYYLiYIKWqlHk0YiELPJO1JSFh
EJziLfIUknN4oUNecGdGQfHNvldO+NgLZE8ysRJhJeg1qwa0GKk9svqIH3Nzfxvl
ul+YgWERCfdwksjeEcTFU47TsFqyOI9WDoVjAzYJD32RQNwSDpRkee9uqyUXbtYK
ID1St/J3PU8SeJH2iNd9muXudx9De6qUe/ppk7o1VqRL8jrZXgNltR9hRhyEH54l
BtzMrroeO0gv+aIpbKsYPr+6sj+f1nqqg8G9GIrV3gmKmTcLmD87LzTugeIcbR/1
OHA2OU2jm4/YdrCX2MHmqzvstee5pctrCF/jhXQh9cFlYiivErxBFtCT38fXGcqV
bWY5gTATIU6OyU8daYFg7e9IOv2D0aPLNmvIsDt5Wje6noorNR1e25ehWvtPPhdO
TgFmyFzgpXPTmYsYvOVO8JzIPz5cSr77JlsovjZaodB6yi/2R+5DjijrzQYQuNlX
Le2p9ruGp1UHhCWONV5ABoHJ9YZSAfEa1st1y1UJoRMqPsaImPTjn+0NSG/NIu9v
waP7Sg14pmSqSa3asfTQguhuWUMYUPZeJcETaQzuYvfAnOf1DRgzbpXXv2uBdjGg
Q/57XawFek4mxgvpVfLqcQssw/QlzzJbcB/hKw3DGbxSNTMigEMxWNNLOdserpxl
G16zJGCrISGH+UZr2HFfE74aCysEjbqOLTIiar+2/08X83RFznV/bDKVmsQ09kfT
Embc8cMx8i6ztqJ3a6mKTRkXalQNCpzPyveHpsbnhw35aB4msSpZSnMLVvoaNgHm
pNUBmmZy6iuGJcqBN+8hqEna/+xSVCzwAd7DzgSw+z0d1dCleDXbsn3i3OYV6Ka/
KXnS9QeXIXxoJ4ivmkGMjYVZ4jjpNCBfjJnK+3BjsmrDFIXcsEfQkF46mJkZi00J
Rp2BA7/8eKFyI3w9oB6lGWAy9h/pws3LcmtFFPgz9pGWxnJXYkAflsOX1YLosJ1+
VjRp+EmR5+aVqidyQm9rOUg0gyemcmVDPi1DA+2FPbla0uzZOaL+QP+InBPuirQX
xAVt631FCU1dOiWBct1R545uX+oF6yDTpQIokf1PhVfR8lCSe38ROYNHnwhIIyLq
3DQVHI6fS8UYnJW2e+SrDouxutbiSZgl1rXA9aOcw5heLoB2Qbzsl3mgrCExSTfV
X7XHaeqkIQFaFkOx+7Qwn/qJgjl5GL7CG48Qwlg7q0jt4JHoeJGgiCQL2OZZtQzi
RWf8YXyg7LzupISyh/6eQpZXmE34bVstg7Px79cHmhrNui5I0I54NryyYwdkIjlG
UusgnQ1jUe1/Zz7EXvgfkVKISJS33qJ/eP+JOQIF/Nm4weo2N0WDJq4jpNKZFBzn
ImYSarQCdSJkXB9E6Ojzz2oXg3ohceWrXuaWZ6VbWELVdJ/AJwlMH++WADf01p7R
eCNz72RAFz14Fv7FEKgEwF5CQ3DIR22BpVpbe6szZ7piF5ROHevUSOckHDy8KAr9
tyXoQ8sFBBrOvHpxgw6UP5eQkOZIj/g4E7n7ZQUcPj22sPHgg6ZAigW1Ij9+Mw6k
NDnRCPmYBCxm1P+mIn1jJlboigTRcTC2QuFqzNvYiMJoiUhiug595JuI/x37AE5i
C0G225b5swGjSlfzg0yF7NBR9LYojJsZUkXFGrulOJ8kllsxocBW+Rw1d5LsNhb0
Qb3Jm7LZ6YJrrxMbWDOLLWpYqbj40hb/Nals+fzrAWGvmeUUgpFkoi9KirxFRk/N
V3EznoFQBEz5aNKpNoZb6w1p5Nk6of90JhvEbLT9gNUzNlR1AuH/p3X5V1AAz+8A
cTHzReNT6nPxCgMRoS7f/7swLM+tUdkeGTSKTfNGnNuLux4ywbmdY0i6mRe0FpmE
z7xTsB/eSVy0iPXs3+eBZ2QHkY60Y9mrX+uL+WKJk2RxG8Sbv/eAGtoo0gOouBVD
BHJgLkkUk2Eg8DYtxD8qt6/oigcfCAulQfRXyYzGR1A844Z7tHv6QKjqUVtJa+X8
T+vNaYrOQBOk5h+cNbX9ohPys5R8PImTMJQjI/ulI8ki2GwrdhgLG7DADvRtX9C+
vCqc+XszR7h9npaVOHfAXYOJ8vLc7Qy9rrHdoQ2erYnHRbiU4nY5sjOrXr8Rl/C9
g6yro60zPuEKZ4XXs7FWPQnUHy1ryyJuSNg2v9REURpuwWh+/862xJE2MUbMhEFd
A82bUUDYKkfB3RSsXtkANgETHHsM61zMHwouX0g1nOmETKYH7qqof1e1TRGvFlDT
vZw5ueGuGwawqrcs27xtH7tXDAM2OhS2F+GvXD0NJjWljX/tPRe4dHPBSbvpaVxM
LYBOfiGnRpleMJ9AgBlFYQwX5PQ4orfpeZUrb44v0LpszkEweUX1ZLLylOUxz6Tj
d8ru4XFG47vrZTrHETLTZIRiAWoqUZftL9Lg5CZoHEyajQB/+pxHfqMQ5ANZpwpk
7KY7eCArvfNng1XquRi8PbLi7GLI6RVyZH2XRYHegVw3X9zJUbW9aY9m6ym3T34F
ATjcobDKP3DbrN9Dj/ECPRGt8AP0HGT7VZRITAch0GjzqqNkkgdLqwLCqwQlF5mi
jH6OJQ1qnoZmk8p5Kdz0jne4nk8Ri06c3Y/UUE9AVwDSfBWkA3AcpOMQnh1kPfO2
0zA42OVe81cfldVgHdZiqQjGpeldJ1AVyqMZ41nJvrCzNMAxRTPkvo17l3TsS/T5
Mu0IV+nta2g9WK5ZDrfHX0a8b7pULdATp8P26jkziW2Mfdcp5jMdXsssNCtrqls1
UPFm4S+mxIo0BHEoTM6VLVnvmBR51VtBmGEBY/1EtihKcHpfBRGDDBAxxFPE3Mjo
myQsQYF8v8Pvc4QxlR/A2fMCy2XzMoc6QlCIniQRdTjadp4nCJ0ipXUtyE6/ft4Z
VGilWsuWB213C3TEFeakQKqLjeTA/KsD7WTj1FDMJ+Bj2zWWDefFHrgQfseDkkS+
iYzk6RozyaTAeQeA5Vas9OxduJy8AESpKRsUfz8uorOM94QlklQ7ayO1VzvYLMWe
G0+xe2jvs8AIwiFzIX9kOIau/J1BDTKXjQ4gB9mGZ5tJHAW7HBAYDLZFL22x26rJ
bfH2MaTNMIYwzfVJKMVmLydeNogmnddMafCg/FlQEhIlLj4tViPjYmZr/db1U8z2
IZJtdyDHkUlHEyZpdPWUuAC5Hl9zurtcU9GA3I+qLoDOUS3q0baPTPsLnspIlOOb
TA20E8wsQsxehRTQ1CVy2ff6RomRlOBtiK5YgkgTfpmVdqTQuzFoPH/qLvap0prq
Dga161xqFCFTOV5u2zQftjvZUvbvc37Mn8uZSVe7CruVJIQT/SnjE5AwQ9skHmkr
F0tlWqJxfZ+S/5lLvXt8VDEUMLz8c53xFXgYeshsX3PtNl/x0Q97PBRShiQr/O4X
/hpigjH++UirVPzCVIw6XAL1lwZ8Buq/0JikKknVjYI/k0k0IFaTh+Fo2IJH7rdl
boIFLnd/EuoyQen0XvBmGsbYMcJh7Y+Atgz3xq9d17i0L/YXRTtPbJglwT4ryyhP
vJdjuJYssMV37HjuPu4MDTjg7R4WXtEvgmBom31Im5Q6UqCQSgmcxhTGDQF6ijlt
EZ2DQucwgI6ByujpJLIhkX8ioZvy+pw8jmyv00hHJGcHcSr2hELJIUsuwF1QY1Rx
Z4e8VP50IrPOWb04t6eWiVBDRiqCxDwyW7IGx1CknY9tPbKoOJYCD+QScwBFUS6M
FcamsHLQtXDDPpoWyGEcxpDiZTHITDVKBjs8wR2VoRmtmiViNji9tgROQRELvRND
BCS3XeM0k8i0E9lx4UEOXQfGA4Xj9FVp/fTOFEyCWAf4LRYII0nJCQ7urQ9oXbOy
KMbc7RhXhB05UdcqDGWquziG9IPSI3bONETcUrao//MwA+Zl35vNI6ZkFONcPju0
07Ye7LG7LBFaXX6FEvPHGd5owGfToM/3rN3nKwhx/y1/wP9WSlVgNDvDUQsj5UEs
DCIpxi14tJZCcdXNiEvbidl86qXakjklT06XPLVwPe51Ey4wF1jjE1qPg8hU5/SY
9ZcX/ig6cmfojDTw4uUAaaq7mIH+bp3TYBlCLJSYyD03nkHAIMtR/IABCwwGWf0h
to+tgORgYlDF55OtsoY9RGN1/XxkU33psvRlJPUwy+QZ4rF3swvgIOKw3FNZC9z2
HDq3+GQk3f+jiY4VEl+ljUb0r/u0kjHPa92n/1NqRYjievhMg3gjjZ8huFzgsNRf
qG6S85oHbrAsWym34IEK0AfF5448uM924/ZNNxa9z2aD3JRbaY4PuQnobPSWreSj
n8TFKFMdEtwAhiXvn8cTOZGq0rJRZTsEjYrfvl0NPa9TPsqc0pe8OOV9HunoobIO
EBHO4PhWYDHO6k0nN+a9q30kX4Azqmor1HOgqdAfCNTGq4bFUpjCiFdcHfkgdiEl
SODMe6UoKvksfPJsNYX8qVzfdLUOWQfmWpjWnAtav6B64NnZhAoONVjrdg2BEzkC
nXkfUle8LrIoL7iiMiWvR/ibBd/rXD7yiAQQVRb0QifF5cyFol2481VLZk2GjjE9
/joeIuLwwCG2G+3g3oCGtXBdGin+NsagXsp7tEi1gLhVJEqaWUQLoQbwdKJ0ECuZ
Kc5T7PNIJzE3WZg11xl0cpfGHV4/IZnQAGCCsb3LZUlVEksiXL+oMkam5buDjrch
P2jhpYjlLOaC6HuE0vtny6wAYb6BtPAfGy5DbaMSjRD5FhaS5B7HWszI6Eoe8MPo
u+ZzvsSROognRCjZE/LKht2qHYBWOjY9vPR4qHTdjHBKweK3bbtzmJ0EjY96b6Ww
GVTlD9IgnWa9KrRcy23BC+F9xL0yVpVrDASzY7JZ4UN+Cb38simWG60qAYfJSN+p
zXgSdHbsQ/NQkCOTGiBXKo5/ztFiWYhS16ScgG+/Sq7Je8L9Tl70+5MQkX3/I/NI
Q1U0HZz8/3b7dklMubwRtyRQpMLvTgnbjKyraGzbaHRA5b9UVcOG/6g/RvS041z/
+OlDM3YkuM1dhpczwEzIN79nMod9CLAzzCoIdRo0UY1CCwPV9AQVX0XWVWoHJ/jd
Fr6R2Xe7kEFPf4MEyFGKvLf2VofnIo6Bot65aemWhyEn3VIcO0yhyWJn5vbSZ0eG
JMIVTuQW0oweFCbY3lTIn/s6S+Ou0iOBXGbutte4qYLSjFL9MWFQAhenfw7xlgEg
Kq57zOFlI2J+f/sSVYuTD1ME+IH+BBkjSRwUAqv4jbs3KtsCl6fjcYLrNK+LUzDu
wT7ispQczktk0OMJgBTuEbMuEa2l3FwYHnxvMinJnGOcxnLqYRUOwQbqxoOuCkd2
9FciRynMA+MLE1ifFG3Ga1iZ7HoExQZYKAAnoTiI4dpJbWdLhiFSUF+cyD1doOm8
HvyCq6ujxzn/Bntq/VMy4UwicpU2i6E/Zd0nISVTuhmEASgeoeoXzxGUb/b3CJjY
JnpQg8gXdXtPonwbMQ+ADofwKRBGIE82ujpWV/H6zbG5FRcj+3JPSIFOkx6C98pK
V5DbRK88G3mwfmcN1QImazIxdc8JYcesqTXAZV5salveM/TMZBX2tG0OfBPbY/o1
`pragma protect end_protected
