// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:54 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
FsnAYIXPxLOdaZsXHqSiuQ/Uqi9rd9+/siE55vJqfCHom35mrCM8kcMDbV1wZ+gC
oIXaWk59LEi8ije7qvb4B7KQiA+W+QE+hXskhBxclWHK7Si0fQ63H/YnoaT2jnHp
oxGrA0VrpGZoLrhiglJt73yHNoJ8+/OwoFOOl55VxpA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3568)
b+SwfRVbGTcaHmbIhc8z/9y5sOQ2Pv42GoG5fur64+odrFdhCpz7zjC2Rf0FxOYM
7ogrYS/7GikHq7VPVpFwkgkjAByFObrhqt6bWYpEawRfmlLcXvb+OExmZ6sGUbam
NTv5GsLhCwCEiGOQG/VVG47kSwglAor3wm1cJgJAkm71KkXcVRAvvVofmkhWZuUo
D7s/A84bhXySkC0MihpXlws2DUTRKdRsyE3gL4GoRrVsiTDJoZHM5CCzPEiy2FVy
TS6kCFuAU82GEqZQvDfaQMKLUoeNATOwSwbr/ehheK2TJmtKGi0M/HcGZDuI1Ocs
ZHPGDtSKAVLQPk45LMvzW05hew3ThZ9Wy3fk+WwndcoPNbyGmh5h5TP45D4iSEdo
mFNZJgzV07zagzwlzlr3JXEn1tUdMI54SZKlWULnEJyzJRcoVtS0R7pJXCUikLG0
9EjqE10b/MPpRDPjHZqayKtpEJFNsdbu5dKyKwUYaEHyOn0EMqSm49syMPRdRIHI
gib5fYimdc//G/DD2w3cThLdjtSWol74veG9fZDXdFPSmIODsDZe50xIIzA5yuSy
HA1RsaDFxZZPMCrHEgBifI6fOMAtgpGe8uRERyair8M5SdTaRnknqDCYX/Qq9tpN
4lfE2TCjB/Jk8Zy8VxuU2neiL+cmCXXy28UmJwXIGNd3XnIi1MPben8NhpYTN7Wp
jOVNk/lagqrozr7I04ZJyTWvnLKP9ecInnJT4ORnJXwcHyYnnuh4pOHEvgK6vWdN
CIB4MokRE6BV7+yIIWn0hsXOGMlPj0fJ6HBRsNF7dJy1wgQXxrOj7oz3HkmAGSlf
5qcfaQuQkgzghDqh9kADgXTJA15Yp15NG67xf5Fegege58Y6dRBO1SzqyiQ0wsX+
rG/so0T3/xE4ljHkaS6TgxkOqPpGGSNHjXvCcj0JHauOjh/OKt+ctZE4D8Bykxv7
T9b21+wpPy9jgM7lM6OoIFpRsd3JN6xfkzG0mCxTyWE9LTtsbQRkoUkmHiMR8gAD
ch8q5FL1rztw1gzrH9eDIAhEjFpSfLG5FuPtHQmns+4O8IF+8gFl6q2EkTDAar6d
p8mctJNM5N9PJ3qRzZMec2EWGDMRhA4ik08Rr4KZwR5+MXA3+Rf01bQ6mqRe6hwt
jLGMrFHpQiDkxydGUkXeiFUfG/VL5AfkrkVPnFxCAS1pxF3olyvLC3lUw4jhDj61
DmDpjzyOT3C7jY+33CawA5H/tRL06QNQQMWbwSzoUOrQEbC4miI89vw6qGZynNye
ptXHFoomPassq401vX2VoNC6I3A0Qju7Z+z7+QPWyWAEtWK/hAxGEkdT21e1DgWi
xUdxQyiE5iLqz3tBaNAn49S8uJCJi9buk7czkHJGxGjs53APF5Cn8gPh2NHdJCsf
ZdIifE/jEOKphzq8LSxAfAEa6hdC4uqYI7r6VVMfHukSg3QauV0+P+cOqD52NXnK
WaQOXdQoOeHogth29vHHvSINhrVb6p60T6mtFmbRPXVHylt6pyLLG9yv7QkX0c5r
ko9ThTtp4f0gP8854Ta8JOnss0FMGlOMW7f5HXlwR3bpZbggue1blXgH3Z98q0eu
m7ajUo9lOsNbghnW8iCuSobecbxEAcrLYFvBjDeHfxNpnReUkyOzQhCHovtwmJyq
14BvbwLXt38FKfdeW12pHCOeKj2bjV00PbEFUReQbZOq+LW5tJvhMcl4JwvE0FMQ
/ex01Lw9IJ5Xe6/nswOdTmVBaZSIn5PvzdH13cpV5i2sSfGzqPdLaCoIctxBuCiX
++uuuh3/kEurvIaTgbrN5iwVcoMcdvzmWBJaGqRa3WwWvj6UNVLh+68pWCudYadU
N3A7Oe2ustFmkggSSZt8llodrbUgTzMXHSeZw2yr0nJZQ6/wz7RlgyIUliC21HOw
pWWggcWbDLxsU1w3Ffh+cIllCzDH+WatXBSiW45sQH6RTePJ2ZOb1i2a4ou5sVcF
uw3ExkrZsj/riQjzyEqvhWoy27IblHgdxCbiIm1LJIhmwUQa0YRicsUi4uJdEQWG
S8Gya8l4EQLA/Ayj1zMLGwGjHeZoVP6sVs2udULxUM7oY2+EbHRBmQ6btY3i5or3
zUEmAgvp14i03jIAGnwbnwydj7bgmB1T69R754vkkhO52tcDUGjz+3Z2rPdRoXB5
lOEoOLZ1n3aH4frJ7Z6i6MzxDCL4wl+yRlLEayleCla/yb/SC8BrENuWpWBVPAUe
xkXVYlYiIgc1Ey00+ODZ/uLZobx7vn2GafFVcibF3cWH/dj1fJxXtEfLFi6MOR2l
drCFmLYTYwTMDK+YTyqv7X4tjuSAWsfG/Rq8AL+zE4TgrTHqmTOICDIyM6DxMK4x
w/+qVGRc1RHyvdn8+mdwRcTs1NwV31d1d+tg7Ysw/XleABM7LyxducTwLu5r6nH+
XOBqijWRzeJhqa8uLMCmAgNWyEmf9FhrnXADd/bGldwZIZbcXzgfWuSQlwCvWTvR
aTpnmTPGDClGm82b2PTm9XZLONdI5ShFIUCz/KkO9E5Z3hBImPx+IsZe5VIUubkq
YmA7ptsWVrzvgyAbo7kWFVkOUuWRDEZjyqLHyTyzBqPb19ajDMtCkdfFsRhfcT6j
8sl5fcdyZQQ3p4EN6w6vT4IV0xLsxAYoLiRL7rGuL43dfOkQjUqKhLwtbFJxqgDL
WuLql/NhcYrGbt7aUurfbHWmfRPwisnEy7Y99LBZrKqrBGAn7blv5A3jTpyUqZ+m
liTgcuFnz9De/RGRjrsjvcVAx0b+zq8rUPat3BOJWazIHZpxZ/1GitdseTa7QzEM
M1y350JDEA3jbsJ5aQkw8KkgAELIUHY+vsHcx8rJxe7LGA3vzpF8yw8KkLIiqSuc
PTeLlSc+H26jhWKxO7etm/7izIuk5KAHzQ9QNRI7zhuEoam8QxzzhxYt8JjoZo+y
P/O1Y5QS4b7DVSrpkpnZIhmjJuNIEV51ZZzdFN90FAgaxJd18zN9fDdXjMAswEiU
dazCPICanpCbnYWzhBRbyh3JRoTGkdnmb8qar8uP5qYGuJGNiJnZqmVxc/RLncCd
geSj0R8PsA85no57zVbfAUkEj5VyYrk3C86+Nc/vRaMKnOAL6P1dQhDsN4B6Pd/H
w9s39iD7kjsKYLOIFlzna6GXgjT/8qOHOLJGu1n3T8TxSF8J0EIlXyQvhm8nAMaz
ZbSngUJVeUi6MEU8cpfURllwXZET3g5LMeAnHBZKr/VmVa+xZLlm0Ex8tHrpjVLo
iAuiP6jiWHOgN5O13PkMmpDMPYPmivWwuzwMXob4cHfQemKCJIc7xe+zx0JIvpVp
JOBOkUGg0PwrB30JO0xjE5OTbJJdYSuQbKHPlbzhI0Sr1KR643ACM3wVM3o6uxkc
m38u01TB1gbR9leUhMCusumH2wMNASnRtc+TvfPH1Zk1tgEsZ8qIJH9XRcbp1PMe
fdq1LROaIBcL2B+RlTcA2w4+wN69KVTnKPZKJ0Yd1kUdc8Tr/xUaDCWW2Uh7CxdT
aG12E8OJbRF90pmIIv1roWJDooH8A1FaNihS7v0eRHsJovtyJnI3hJYVdF7EfIMU
9AFAFxAOtgqCoM2+E/9st3tjpNWF74lfCJcYIW8nnCF/dP104qe6vLqZNccLzOPJ
jvRi4BpmsMZOQtnArmxGsBIUHtAa1I5iK7RgXztAyGn2RNBEcbt4Ek9rFZgKUPZT
JpyC2vMIWakssa+ELbX9INX6jb+7JXM/tYSiWb7h7LyBlKBpqPlw4QkDIbQucbyS
G16EQtnIpgSldnwI//JXbL77WwOokrqCGChRi/5b8cqQUc6bRvgUfpIL14ESNF+/
STwRykGaS/WymJunylmfUWsjaw3N92C/A0zWIIXuwSgH9npNFKFYRT6AwGov34cW
0yqGkCoE7eo+QC36087Pnlks5gtXLlBiCkQJvAz+p1WpvMuNt6EdEXHNPpFM4A9n
Siojle29Ov20tEYy1o7C+v2V8in3N0HqHfLB704y0V8W0pm7WsehociYhZdpdDOM
4ZShotD/VBtXVkw1evIBbpENw92eeEnzlS3+JaFM5YmIWu5sjpeZ1Zaird0cDHIz
Q98eNssNMm/J9IrZerG+0tmRObH9RG6hWH4N6GL8pT2qt6ryG/gAY2U2cL0RA6g4
sZsCV9JCP2hEhnD0Sf3M5MDpj1VwPsmLbKqOkJ7gpUZjMCxGvbVw7cAYQ6uTVB8T
RqcYlA02rfWbvLqAFceW8kylCHxlTO5uA23J04QMT9shl6Yb7kygFnTPJ5B8psGE
8U3bjgl95Yxxt6g61pOpuWOYRQhQwKh69+W7LwyYVOjSOahh2VGJadAShE1PArmU
t6JDREvgKWtkFUI50j3JpyHkIg/Kzy2PC5gq8DQZpiZMHBIoc5cnRZZTJY08HtxB
LW5YO46KcF+QeYQ+YdZyPbqBCFfykvPjnDLXfueyWNqBchT8ZzAnEFtd6X//Ek56
soLPx5vqC3qahXtc1Lywv5PbSOihf1gCAaLvS0KQZcTry3jK9awjtTQu/k0h/4b0
E3NCPnvq7P5yiu6pd6Rr0G8lkYDhQV3Voobl7BAgsRUU3+MN2upgnM8XBue71wwD
j6RE7PaNlT7oUjpm8AmHZzP7q3aYC1JnRV7G8/wroUPCVsaYTEmX520NII2GcBHu
jUUYJ8/MJPAwZDRNf0xHSOwBGKhEDJS/I6h9O1AroNVgwKqhn2tXEHF5dPEiFNsU
Csk7GReGu3L64LAJo2EArw==
`pragma protect end_protected
