// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:51 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
WNBbMZd6RQsQGm0kIMkitJQxyQJ2g4Q2I4yZeEGFTWJBr5bIujqMlF0tR3ga0y0b
GGtd70AmN7yLvoMC8b04L0/jg0M+ywbMnl8EhvqblcdDThjxXwrfBR/I9B5RYB7r
COOjO5dbinf9ZjKFiyUxpPww9mAZuepW1Iv6GI2Dpio=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8656)
SjTXAYgUssZ8454rDTXrTjO13h2uWZkByomt2hWZFS3AsVv2v+CmElKgoAh9w+TQ
9enmLarc+VeRy1xBOnRpHe6Zu7pV04yK9o5FVYSnGxiGXJa7pHTTSZYih4uDGKYg
GaUgxS2jTRqoAAjgXarHkUgWDVmZexMDR5RFR+mU5AUJZQLBlPQSJj2OCwq3VqIZ
kn5wrUvy8YHPhuXKxQ43gE3fqpGDzyyKxWUCRSd/8cWss8XgvlUc2lyJmC6r5XAr
0CiVdU5ig0Jlzo3w7ZlVmvH4ExVcA9se7FhSep8GUhP0oNWw6wTk/SKNxLl2fiMu
R97DsauZGn7223EHdM0ue6whFoZoDIklBO6d0Hv0kmxxwddllfxKCMSb9rkMa0oY
kVMpNNfZwRBgkYz/amEhdhtQLh5ufKrJpAoxE9NgLc7w/ZsVf3yvhA0yeQ6ZG7TQ
sapBDhFvCNM69rnj9/WFqdd95W//w2eTAYpURRI6N2QvMvqidfepwBAvVa9eNklD
B/ZtTwcePYu4vt/Mr0nqjBmJp8OKryrap5cAtJilLvnnJ8KDaYS4wD4Q76XD4v6g
vvVjaWuu4yvfcELXKOTRpQZ0r7w/dXvgWgF1TKjSlP/+QI9AFr0YKOXoGGs3LwBv
yS9nPGqPoCeMxvB9wM15uzPg0f7+SZgBhLWu+nK4BTlhFGUBJG+vZZxcrVgOB2o5
4do2yJVLeUZyboJU61fbxp5YqE5XWhEPWICKhY8gzczUcdmorSzJK1IVu7iaEl2f
yFU/o4o4TGJmSFcverzy/5q0cjwv7F9gANGRNi6zRGi56B+cVEQRHMCc4PuOF0MT
WpxMaBHJkEsUm6be3QZ+PeBrRTRu1bbv3vqh733Br3TdNEFU3h+o+RWfSnxEYLtU
vcx0SGvsqa1FNqIYsfoeowoqxeULq76pkmuFYY4A9/o+0/BpIhn/gUhedrz64Tf+
jz4nrbt0hm47x9mXxP4pk7Le/7+svKoz7f/kigJXB7Ex5RlAfY7A5asGW+3hA5sC
1r3ory05VBzVZFWA7bDtNW86NGv5/rRgeVyoS2Pbg7DR4psvUUw6XxQPjVtNC/HB
5AqnR7A+8qt1PYiviAQ3Xfr9uBYjH6M70k5slyby8A7qMw3QyGNH3NhPoZYwFQVT
TkpU5CASpgW5ZEhXQcNcy7ZSRwFMxeXkYgBvrWP4L8W8qtNLv99oz96IwvzEZ29j
klMddc424lCI67h3i2BzEWR/pUQJ/tHFfGnENwWUQhJg+njDn1EiftwUG7ab1IFV
8jNNh4/MfSlzLrQZiB91NyDiDBr6uehNC8f/UtVtlET/BF7EsH81uoGPUhuUMs3J
bp7PpzHLdGRr7FwEXPoHpBtJ+mPA4OYfyJ2h7N4HcZwoX7QoPsiYHimVrxtKX77l
jB649uRUGZCnjItYPP1tVx009hJEvodeOZRkcqyrhJlHcjcezd1VHqYUXnvLD+IF
OXqpeeTHlbCD/v+gsv4FD6pZJRwPpuqQPowgIb7zGFU9WR4FvK+Yv81s27I79kyq
j+om0P+VDOGbVe+Q31HjAxqdZkNZhICxYey/Ky3WAZHyZG8z3xToL/BXQ0AHyYSg
0a9cpSokmTWx9k2KSiKttHI8ho3gKxIJ0SkfDFqE9IezvpYuo4Kwbl6RKuWRNNDE
5PD4g/KzpOqrm6K++tJugGLtsd7Gyf2dOtXkkbI5+jgnBcZ/k1wjEQuXexXw3YKM
m5DOX2Wxo559CVQdX9A9Jfwmx5EFtwM0FgxAh9a+w5x5nyTSoEn+f67lHAcREElI
HpqZmWmoNoSkbbM38hNv/5vL7aL9xDA7bQ+7zwaRLRwqLKgjh/0Qkrreyla5MgsP
TY0ZTRQaFjTrIzuH+m0KXW3x5Dw0f2qL1xtnLpWx+ZJMXKsQyq533p5TfGb4pP+V
VBzVULQR+g6nPput+s/VcBosm8BHXcsvIHYk2wwbdJQI4vsADuFWoRN1AO8z0JmA
Zfb/rQSaRXLs+KLbCirKaQxjnV3fGoHaJBlCXbi32StCQogcLq9F6DC40oMjkH5u
FfaNOcLqPmBjAiRyVGX/AKiG6L7JAAyh0buchGrJ2mK+ZYK1hztclXe0Iii3CVYn
fHcT3f2JGKY5j8shUFxTB3yI95QkKl8DlhVzrTDSKrRWaRwCgQWF7awnrU/uaxRT
VDKCN+wI+lFKt2WaR9KI2F+sfoSmNaTEsPpmpYJMP5Ce9D40RyMOCBLH5rpwV31d
wJEAOHtmouGPlNwPRFh27S6ZXwyW5T8SMiuOgU2XvVxs6bQceyV0UbTc9XXpglmx
qbC8BF59UTxhVJPBDpEr6UAf9w5lD5lipbnw45UhKP9U4Cy2+7cL/TMd6V3Fmvyg
T8E9KhKgt5drYnZZfbbGjKd4OCtKbSeMW10LqN54oLImdAgvpH1tujyDRb7pp49g
K/0DC4i68EO/jWUDqDJFNTLVoYtRxcEDpu0XUO+4bQ2V5IhUlI0oP4HbjN0xp7GS
02mpYV6jXg2MlzLQBK8bOxnFOM66Z3aQqmaOklYZ0NTrBqubOKsmgKVJVnsVut1w
ksCYhvv7rNl3SsO/LxuFS1LhU7MhzPgxlGZBfcZBVvD0iRR6OYx24bnpEdeIA55M
0w+L+D09khSsS5xkpxGyZvBBXfBFjg/X8v/lA3TsOh+BJRsL6voOex4A147Fky/O
2KQhaC7QtNQXwIrY4DDhb/w3Jdym7UIscuqmAU608UvF20pkf/loolr8UflGL8Wa
KfXuOrXat4ipBIdaMgergZ6x2naZmZlNgehC/OTKiRHgMp93/8TDevPN0dQtfAsu
Plo0eg3Cmz9S98pkMLB+9InPnbo0YPL9gm93suL+tPliLC8gKWRRBZaW6QBP7kTf
tgiiKEvsBCdXxdrUr5n336Lp8uWt9Hb1CMIXE9WYlo9cLChNvuk5eTR9V752swbG
OMJWju1NltJ0L0BcwM5eGL5RU8yaRoN45+36AUjFRwxSYDOp01b6KCBqozATtMvn
sVZIv6DALOx+uuumWFeG1hHE+UGQadGcTpa3sQHQhTJQqbUEeZiMTA9wC71GZuTC
wq4d+b9dOI0E+Cti7ck7y3utjNMN5VrYA1DzpbKo4lC/7MlNT7sebl3EyvjTvn90
yf/dsfGcYc+shM+N8fouzAF4Mom9+A/GqHDsuxcpw5zhUF2+r0RcL3X/xb+jW3FV
AMP4TPYF3UMcY84Z8OUK6LqPtczLfN4SXjJBnCRrfGEoOhQOupr4BYFJipRkaz69
jz7D2VIqF8iNeXKchyh5DEreUwLdYuUHI4VMto3M3a3+5Pc22+7RUVE7HUsmCOCK
QaNXo/Q3Z0ENSB9CjOH51rF13jWHJnFoYeAvoJwCSRXx4vulE9ZrXw1wfkGZHvuK
7Fu/Yv1AeTUmM/wKCpO+ITWi0ZL6zeoaDpC5CxNT02QOI8dYxCOkLQum4Ro5LICL
+uhbiJO6a7P7OgsVicLGvOqd6wgcDZ3w/N2hNF5yAWGkyjbur71/iGqhFbHSY3tR
Si5cYTosfqTa8SBglujX9FJTOWhHb6X66U3Z0tlsxMfWwsy5WCz3Tgo9Fsi5PtuK
Lkmmjb62dZgk64vvIC+Ztn4kHdYX6wPqs//oGjfaCySJj2N+wYlSynALbLr7hTjx
8U0QInKZR4h8VSAQj/tvXF2YvOxyicCldp7VGzEGvPcggkuOxneuvO5j0IzX3F7L
m6HlTWb1MXAcxN6HhDc+X23RzCYVW6etMBi8D/Mnec6JLpd5b2gzEEdh8VVzccxB
xQmbwYulI9wtqFmzv/rn7vl8skGr6M1+oSPhtyJaO8pNIAiyJ7A27xWWSQROj1EX
fklmlMqv5kWSLLxWoIVGlkkn/5np3TJl9aSLdkc27N+EzXU83/52PA6sbzL+cph7
vjAI0MvWMrS6QrgQEYDTm6q8K43Ol5bEID1hDjkDDScC/psjwOnYMWs/sw5PIs63
Y1pyp02p30Sy+0HQlus6eyFXovnJ5rwGVrBw1io17RpaBYa0qZmGyw8R1kE19lny
ZFHer+E4eCtQwURdhtVDcWR3Vji5m/vKV3mXyWJWO9tp6v3N2j7tcbaq2pCiDtNX
bWs0OCXNyPP/29H3IelH6a1HNMAPMAeEKXoDveKdrAx18UMGJRd8HB7qJujF9gTa
WfqCY2TU7owoU25PN9AWA+3nTM8/K/TGVKfSZX40WWN0oN1IY5+iTQaniBWX+jHe
R9Ce3gJpgMXrchguqvzAnWpSgZ+MlCtg2148lndpf43bmpJFRyOfNdDdI2SyAsK6
2vKt325N7D1nJIaLB1hqy6h9TPeDdXwo+Q9nLGogsViURkYGsUfjd8SFdUnFYbBC
xMujq52MXRJQtBo7cXp22xLc4NtUtcyFU6h+3gkWp9V/34P75bYSswlT32HmNswb
eAEkLRMV1OHE8dFfFfvqJPtv19I+2wMuadx6G6rCeq3DZFP26FwDx8nJVfQo0Wg8
6q75FhS2PCwaanCqD8OqMUEPttlLoBV63Fdqy9hdEkKvFpg04qmp92QWO0r97+5r
PcsSPPeZYkcRvDLawbUNMlUKmqJyqES5NLMZrlvgnbeiorlF9N4kXi3DjW1Czk86
DxwrJUl9V24/kBV9RpsHEo+UKGTKpKiYP4sw977ronzX/biTG5b/cEi6hLMjpybp
lA8SV2QS1w+fO+9GgsNZTXLw+hwjx4NY5WzPDWXsQzUJSAdiRCI1SixQNxxKigCx
vf8ny3mobYMvZH+qWLrA0STTEM6R4ON0R9curxYdWoal85kjgZ+lLqtBBqPxqayd
VUcpg8FzBb8CSL0LXcqGs1iKPv10F7ZKYsDqWuYB+2sFXwqbInYalJljVeSgg0fy
uSlcCa5oa/+Rni0XdQYT4aKCTjqjVkfeMU7QvrpTi57fA/E43q+0KTUkbQ9ue2hW
sC8CiAHIWT9ijeaNn84VAPzbz96hhaO2LerWeAHfEjJdHt2A1NP/xaBZkcgans/O
LPHuNou5XxRAS0rBrMS02j+uS1obDKMYkpofvfXFv/xbU+DD+qYUwNKQi4GVLTHj
QC9IIiE1qoT+n3g5OTbaZYZ/VCT5T+6gMObejNzfWNwfY6PvP7q9vop24g0nKW94
R0SjyIArWLXBHqQknHHqYOdBQjjTTJO1KzDV+PzV+0+WUntKN1/+L6w6Zl0EAipD
Jc5eAXX81Xql3+O1Nou0+Tqi/xKAzHYOmzKtHN5i+CskpNUvit0CXolEg+WUaN5f
ZHdVX+zORkMWKTB0d38YjgOTQ7zY6pqCyXhjsFP2pDpvCpI5Iji71e/CmncBf9mj
lvBVPv+jspwLsI63WhhETRAON0j7ghmRIKloBJjEaxkt9XpIsxg8egL9Z/Z3Ojgc
+9ufsrTJUsI2fhgejkSv/P1d3OlEQPNAjltoAHRqHnnGiF+3ezyQRAJJPOKsY71v
VmbIfole6omK5dkJWVsJ7uIpiBBZKC00RFyepGCBwQQ84GlyQsCksIezBHQQ+9zP
1j560ysudB3CjKCvDED8pim6fkRiukl+0m4jLz37GhdUAjPjHWQwhB1/T2eL/I6H
ZD2UiyfXF5WphpYo2zzyZXv5CfYj5PLlLpV2ddW/vpyakXOKMwpSCT1yvxPhfOLC
8Efa9HECeToJzOB+QQqXjXkAgFctqkKYUhG/YNgA/c6xlA2DqYYxYuiNUU35ROeC
sPYwG7yjlFAjl+tmlPUCBHxEDyQVlzLAR9dIJisJoSLYDrwukC7nDQeLO//6Yd+n
l35jKQDmTjxdy+wz2KsCT5K2m0Qx+BvXPGT/fx4MhrObu14/lAE4YUC7fuEPuoda
Owumfi5bEjNiLOUEy3MctGGT9UZkP1YOZcPEUxwG3QfEcxXRZu1ux1Jby38O9qQn
znq6tEz4Hy4EzaHudTVEiLbrAd4eXPod/f76PpaVOtWOHo8WGh/waFPcShXRvls8
fxgNCafEXYaBf7xis+17ZdbEmRU6rpamjgcb8lYX77kLs5t3ou11SQiyOV0wGo/+
98Sa9Wv49t5Spd0XzxFsCyJJjEhB9Vhq7nSTauCrbd3/gFy0FAPTurQywIYFkGbb
TbDEUllABU52LHSKzU0mk1VhPAGdCq/CYdpkKyrv7ii1xm1V6ROHB3QqupzIHR3y
AhUCgqjzdHoSz/7MaD3akmgqXepI7XokkK7JCEQuYZO9exgii5Gh2TSc0w3q8h9x
ZQUZedGdwiTZZWHPY1totoQB7NB3GxvejOXjQzANQ33nXO34X2vzvIOtbXy1TyAz
CJgCihOgoIHb4ylEt4SC4rhNN+26FvXovQ7KBomwW2s0KNxKZ61/aVv21iaxuBZ6
iw+/rmh5eCcw+/DhfotTvssN58iC5E0fL687tOxi3SRQhxnzzklHXq0/YPLzquw+
c/2tilN/B3i+jrcF50UNSoOHH5bgmL/j++Trmz1mb6gyfT3SiB3hSAkaSbCwhvo3
w+pDetPfg9UdT/Kku2Xu8ZwQpBl70RWWCGtLfYZ6tYdK8UKKAHb2Hr/zbyj01Ebl
eBBNwVMzg626HvzndntPNCLa7M2lJd7WKh5hYk7mfwlLw4cGWYjSYxuWQTtbB2iB
hW9w8Fb0WO3rziM7r03SFzTnFqcK+HpGfIYYuoxoA2e/NG9P3+5CguXn4RhV9zAZ
cgIcFJQNzhSeTQb2YWDvCempISt/RdKF2vMWn/FSpI95robA0WBPywy0hqJX57YO
XFfy7yyirXyghllExnhp3Hqwy/8dnWiW02QLD4Wbmyge3Y1QUm+jolsnhBypuMb8
hx/rssqqUoIixrpVhf/ua6yldPjiRvBZTeBbi2bSnguHgus1zEoaMIO8IEtkzW3A
aQji7YANIi/xwf0Jwa0dorwP9gAywFrzVhgq6jiUh9Assp/SNf9AyrMo4E8px5H5
+euCpm4pvRsGKauaznRJ/QR8/VBR21GOfb3dqDV99G/WqnzX52zBtGFaO2PXv4Tp
FqxBN5BIjt0r5gyeP+Oipc4/dKs9FEffYK/2ihbttpzzrGs8TQaREig/nWBeAL6z
cqno522jnazlrvdK146BPLP0CU7Y7T4LukZhrere34+EwC6KMB5q9KHYdDvjG+eG
m8FURYO4mQaXnYWR4iPIpomUuVldnHdjLH0jMKhU9cWgG1iUVae0fplceZ4HN+gG
sYl7gPXsGnwja/dghiTGofaVVK5rf6n/JINrqHGwGVJUW9u4WYCRNyKoARdNt1U8
h9VYFyJG7AH4R2x+941OlU7rvVzhIfYd3rIbij0G0oqBS7gyATJqDWeXFXNUqR+D
8H/5KtVPTva4Buk0k5NvO3lm5t/h84qAxaGcBjOP9G3kJ0mmroiJ9wD5csVimAu5
6GJN00+j+d62PC2oMechPoploxvjKKbnB8jIbia7/a5VDPjW35fHBh8yd8T7rWCn
WrytzNQdgzR0ywlSRpxlezZYS9MJuiJw2mmgM6keqc/RrqYcJ4jQEWQV5JvfCQ5N
AYe+cR6/DxniUb/j7U2E8J7ZJeH7NUu9jLtbFdJLz3ZGSNzg3+LuX9IYlh7FLWdn
w/KD+4+51gDKx2hieQrGtO2qLNgTjYkoYDtydgGyxfgxjZGVH01Rs7Iul7HqGKPT
+hMc0HgkLPTQi+baQlFypeSQkSbeOciqs4Vg11Ke8K8IC8++JPYmH+1U9mFoHZbp
iNRVVlAlqX3qzW0/j07VP3udHgK9GX1Vb8NEb4ZGaq8b1o/OS3ESil1DFiTvkhoL
Zi7EQv3mhrrp2oy1jSYQgM96F7Bw2EgBHDTGoZVDyCGt1jacNR4Mu7gYTpGZW+Jw
F3jzooTTM2W+fM7MWiOhq4Gd478AaZbkdooVLGiZmMFymjlCOui2CJASxVoRBeLo
IpCNVkj4ig+Ar2C83k2RHmIcjhLMM00W9o+TT7oo37UK8RLThcy66pJff/Q+yIdR
w6I7nLkCdOGXgXROuAiCYF3IwlFvFlSbYvDq8irVWasbpbOgN7Iomlr/NaB3EcWA
cCICUK3lzpL3GBljSl8sDHzf+noUlQD5//iooQbRDThPvwCRYCOcB/rVAhow/8YY
XEK7WNBVNTWDZrZsxxIW9qenlK0hvYWmQ6VBmln6pqqi1LRO6mGlbObK/Qil3sxp
Rw3yPx/qpEa/jEsEaQF5JH+ZwvMMeeH6gWNKqecNeB+PGRbXK7LwzVOgF7Ymg5YQ
IdzdWIwxk23La2ZSiK8q/1DBvCtEDr8PiT/JE5SCDUMytQkJOWe38xcy2/TMx2kL
tIzZc/THzLbQjh1A3ME0RuVDI/uc7YR8Lt/BaCSBSheY7K7sMPbam1k0mHjzbM6i
0z+W8RmbVTtWJQWzMmhwwysXnxv3LabN6zwaUpRIndUEIa5re2mv48tOU8VVAwwD
Iz7xNT4oalYz1jQBeEirzHJPeBaglgL9PLovRHv8uzkQiJRuqIZejKZcZxM0ztNC
BGvOSiRsz2R9KDDaSDL4UbPJJA+gJaM1LqtlTiKEEI6aNPPkRCG3etEy84nKdQJs
QbuZBaYf1wfr5BWqsu1BzJaPIcvAyFN0BnYqEpyqSJVkdZq7gP2HpRQgt/6ItdZI
/z9M9OnW01JGgNBX/9o282w98WRAoc3ewMC8rdTHyCU6/2Aoa0sVovqi8yBs5OUn
NSV3OxQlsPbG6PxB+xo21gXgBuN4wW9VHiQtqnVlDYxJ38NPWMaPNgV0mRAP431Y
7zw8UnW19MREKyRq1FmCkzNKc37r/msHcHxK60RS2yU6BDOtgghK/zxecgfdnNsU
/897y5H/QbNDxRYwLX1C+HVA0dl8oswfGYU3MMeH+KmGaXSNuEinFOSdPtkWKoVs
KvbOLsDpaNqi1kIxFytQ989St3CZIH6R8xezQDeM1z6Qsi6PjMcixoJKGbI1y+uT
WtqxNTz80E6R+EnUOOwOztR2xhxRUN/mBrcTKNWpe/tABiV/QS1vsKIkz6A8oCaC
AtetSsIO6710KoeC5GOH2blT/P/8cacUWqaQ+2KVio/xiCxO7owNq6PyY+gS+Gyy
WjcFchulJXoaReK3kiEyyVs/B5d++e7wX9+QZeMLWTAhcaeJr51mdiThEAOj3DyC
R7kPcD+QELH0uOkNvjQ9A6Fo/BEFQj870mlM4aU+LZchrMIQhzByHfdqspIL9OwH
YJVHeD8wbY0S8tZZVYP43A7WWfTqMfdlZvCoRnUVPbzwt0KBYfk29X4Nv42TMVpm
OtWnm9hC55jRWgZNW6iGv4FvO/gnmY4UkgxRlG2w7AEI5fVGqph9YajnJFXND369
AvZYncVCyoS3CrQ/zwG/GEyuIaq1arA+L6vzZCSicRdqaDqDhQOSAX4InXYtPolS
jUeimMFRJlh9pl/cq1yvxiEiV2glh9SRVueuwS6l4mbZHNib4VFJDpzyZLyoIAWM
p8gF5Q9RVUV4KOuTRyRHWSLdPd4HTQOWPkMQplfB9OnD0BxyVJZPsmXRBFgea+mr
9GREdV1ON/Zycq2G9v+o2xutNjfGuqJBq8UwQXiLEl6gsAGK1HobBJwtOp7LVDkE
Az+ua1G1cRKrT5j4nNwNtkqYAFS0URLfFr8zcq2Mgnig3Io7zhuJtaOn9aLFXP7e
92A9JlXAxIqOMVrv9inBYCjTbK2r3dRsIIrGC2bZAaqeffN5fxoE/WloJThDguR5
aIQHKJ99V/Y8GHF8adkSekT2hr+5b7gP2i6vElunxL6o1Z/X0SlKAuH5hGlL61UA
r5CbISVHV1ElND3oPovwaxDisrlhRykKwYMjAOLXMqhOBO30uMS0LZa7dDxHWEBx
pkjPvEsxkj9pmyTJRwivJfhOCPz6ee8PYeczyZCJzDnB1FK37akwjKiDHbgJXAoy
UjRSu1wwVS/tkeJFDEhsUKKczvQ2oN3xrTsPDK8SxoL8bk1Ryg3XgXv0yCf3Jt68
mr486YnusR6i7CpnFsERl0bNb9ZMaZN9AP3PxyyHGPm/EIcoScRy8XxoFus4mQ2W
7SbDOdq+nmGTkLd3ZM+yULBuyWTjzYe9Lb8fttKgQA3d0V6qvw4ReLBQsNp8Rm1L
C7xskr5k24HO0KZDAhCSdtGqKoT8aRVxe/q2oEVpMZwu3dsZZ1PPzB5mXVRLG1hJ
/LN0SJnc6hduE/Wtw8P47YTBi9dBB4jfzAo06KDCsInWmO7c6I7KfTQVTP8ts48i
HQj+/aVI4A+AtdA+7TmvJb+xUnjLCGuBxZgwieye7u6/0ZQXSGYTs/tFunEKkNpk
qiBo927rjqkpgvI4+6aC7BDb6BcJyGZCuubyywvSqr+lC+PUmvcRFye6g7YUgiFK
6UlKO7x0JjpBR/qY0+OiWqH2oU88+iZpcDKlRppBfHga83P9h1aFRWn68dLWMr/I
t52BUd3Qjr1WV0XAk5i3KYkYVnlSQxdE1LZkkMsqCwZa9Ow4/4+HOUSFdpmWSjXL
jazUhNTMvpuSZdXRLwiqk4SFfKU/WDq3eI07bKddGFEurYJd+CPACfoPKG+sP64+
os9l15aXzX62H3ZJ5NzkHwQXVHpJwS5ZjjZT75TB+IbkcqUes3lPREVDwX+GgURe
ylwC37Uc7mH4KkqOECTcvE4kiK+fWV2JsCEGFFL8aityGAcfDwYsrvjNLTZJTYfR
c/6S2EfvnPqykSN+N53EaMVd5e9Cd2VyYQ/WdlpKEjjpyVPz+9Y1Y+bjO2psbaU3
HEAxwNfKBckTsiKVxetNNs9Kyxw/Gp+nkwcFF/VtABBo/LYUU3BCpikjm9pe4A71
v9f1UEjJCseVL6vXJ/Ddw307HtbJmMhkREbMrynrfZ4SiVpKwCGXBO2aWOMU+muw
I7JGR4IbBenBe797vLBKn4gAnNiPRwgL4NDXQ22TaWcatUgSYALokDvzKIF56TVm
Q1YM62el7NsHkcCGAUtFxZxwK1VhNq8gJiZffr7OrCPQ/tY9Mo9RyvgvTS+K4ZSZ
8A/7QTAlFGBXq1gcbqjHImnd3Ou6lekGLoTVTNzgnz85/aj99ezDuvZPJVzaZcSa
ZehXE9fvPKYscV1ypB0fm8HdpCxxxNjctVu/nHFzd+f5mcGkwyVa3ptMoDwsD/IZ
IsUcbem7jjetNifFXiOf8wugzKvbPk2v0en3NDKFVQpT3x6HJLtM63+CGXuUlHsE
0Br7+YeI+Hzk2QIZQK9T72e0T1B7kJw0vAsixpdcrL1wAp9oeD5Wf66sSDfC5YXZ
CQRlFtpgINRA0rTBtOBlVkWLRI8u7vTYqdgDLwHGyEJV/FCymla8VOUuQfdiB22J
r21H9grloLZCgotxXZkrFJ4XYsnGkZph+bwmcouFejLxTIKsEgRo47LrWUullBJk
Sq5nrO0Op0Km1c7b0ClB/bu1+rlSjPlkJLnhZRzPWy1xJ0+Txn1GcGFqGH+WLmdU
0bP3DND7KLW9fJmDREelAa1uN9RnFMVAlpIRX+ks8WiuwsMcReCsrLZAXTVlq33k
V7lCtQzZUu7Tl/oGVuW2ghNrC9sSiHLTJjbdW+N8bKIIFGV0SEmCrOEtxr2tzcaP
pVk+YVs6uyCYT2eqCMfw2Q==
`pragma protect end_protected
