// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:57 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
fJg5ttER2JfyreitJ12x3SV8AotQbkTzY1KVVtZ7+GFNzQVrhmg8Loka6oweyVyw
DcA74VmK7+UESRHoXndIrmLMOHlC6uwBpfsXttBGSIt7eRcGP4WIJLlLGis/OAEE
j0MPxAhngTm64DhXAxQ0mfgNSCvdcAZ912/cTxxCmL0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3792)
Qn0cXlESRdHNEnGUL/BxbTWrpt0X8pjt9bBdtAUps2gf4U3Fbfc0t1M9GC4mXw4t
vdeWmIRMSdacwGw6NsS6YQ9BS/XqWuimxqGmzKYvvl3RzLvgen1wQ20GQLtDTDGa
6i5Gr7r0wMhwNe/vbcwQfnAPyrQ2L5zOVt4PbHc+ZoiU5CZultQ1qL2wrqMb0Q/6
qu8YVcb55/Q+oQgrVT95sugBUmuhYXug/SJbsJgoFMTuI8Y5Wm9sxycT1lD8cngI
FbjBKaC0u6dI6vOgArWdC4DiMUuEmYcz6FyNssucq8hBOXgEaLn8HDERRCIh8pKj
xFYYaRI4WzRI4s32kZH0IPvehDEuhgkFKlH/2ptXaj3lH9AcKh88m78fkD/HF8Db
1OaBvr3jb5E8wSeOo+O4Egwp9m15tse9FIqVEjd3fpagqyk+NNyI0ZzAd083Z/T4
NFjMXUtgii1EdwaG2Xc64S0/YMpmisg+bnOrRAtTUrOPRanRbhL60ILKwo4tc+uO
j0aQT216e91wGtSPC2Ai/2vtaaqSr1NZxx2wGPDLM37UahECxth6cJS0mGUuJXAp
17EeMkfkD+XBXG/ainUJ9iYeB57yTEkuiOrsi+badH3ZsB9mvOwgXD7GDrkrgdZp
XsXwbC/mmZS5LtGX7XzWM+duv8AI8UwvH9yCBRaYvo3hM5RtNKsvHNDgSA8HYQkK
xYYFx8V32FJiewsCH9DaqdHutuJXDGKpWooLxfItdfrG2TycD4gigfCNj5XcZpGZ
fB4HFq1pTe7g9BcJdsZ2A+X4fcLRGCQFOWVd7+1cgQ0P7SJc4jrTVjSbtQyGTY1d
LPdgpuQ1JA2FJ8vxQiqMQ1RL/ffPiCvBvp0RwsyM7E1bqKhWUniV97SToB06k71N
xUYj3b5OVyH65phPd9z0C/oDL/wC5e0Ff9H9e8fMyPs8GXU1PQFOf3fIusHxoXLL
NhMlHhsNeHlQIjjMmmxBBHw9zPC53gy9vKbExB96CNg8nWiANH9wT2llXBLnax/T
RU1wLeH/2RrjWcV9LI1H920VP2OpXBzbCluC2l2NKNfHGFNZYHm0qPVDTbMaHVsx
5C9TeB1h5eumWqhpnjlNqjVriql+w2TmSkajyNdw4dp4SUs1ScOkd1I4WUHWrF3B
MnfJM8dAyGfsuGQsu/QhX0WQo9pri93tCuSidIyCmkUGdpNHvyNt7E+KbxKmxA1L
2A6HEQ/MjhVI1ucqbFp3xVy84Jr3dA5x4Q6rtVnumzOegkeW3h9gEyO67sLJuPR5
sFugFCE634moC2yzkhi3evVAhPv1/Phk5IlI9ns8z6TmEKkG9H1r4FhneM8+9nWX
isb5hvEGt20aASQVJNSfffTQngIWTHRQUhNyUnpaT0uFYh4VaA+1GaEScR5Kf0eh
bHOHjwSmpV4AqjuY0YE3vrFeoObcFRSaBSrD/CENqOzJOL5jJJ4LH2NFfqMUGXJ8
ww/Su8yM4y6PjcPwlmgAcM1BHraCZXQ4hl59jJRUApugfJA73JUV/S/urNepseC4
fWsVKOn1tTfNUfg3411iogW2OnbjN6oc4WtJlOGEoXLmgh9jzDIzA3mvrj4sidd7
7EFI+5yHhGzNwKrMXUUm8rjAi3AAHagop4Nz+/nIPmDbU9kLr7vXLtIdSPkB50wQ
vAjBSqgzPFyv+uiK5QOcELlb+MZ78FRsYSra3VdAY6IAL8OOkoXPjujPuA8ttmBZ
NKZrrPCphkfjTyMYOTQjtIIMcuwdp7JKrWTK7ijWOD7pgcsD0ytYOERNcE04hBqC
szYkXC6kyykRvd/aAI/ibxmewjD0cgk7FouTWfWDVdmFJoThtS8IjnWkiGLCWBgn
RxYTQRqfQDgSEjR0d9BGu4X6Q+ye2VfVmPk83vqp6Q+hQZOfu/7ZlMmnMfMk//U9
ADxmWBA6mSAfKysmh0SzbRB0kx9y3iwn1jtx0Nt+fiNKm3MNua1Y1GBm+pxwO337
wtOnb5U0cy0hA5u4HkWfly4NEKgKsEwkZd6JRLyY/KLocj3KBgcR4z+sERlUtaj2
oQ00VSBeLUbSUuMLUYwXIZpr2L+R+jufmivyxOfMvXx7dtYk2j6+oDbaM6a5kuuU
z3foTSWEw1GhYZzlVC1L5XyEUDOglKIuAKVl0N2Rul2oMuHOmb0XQiQsgjmx8HSm
T3fNIZ5/W4uO8UL97mMrxkNQZ3FZE6egFNjiMT9nSZ0jLGItV2JfFfiSNjOPKgE3
AEHi64waH75ERFODwhy/5msofwgFO9QR8PD2gBragH52Hr3xVv/oN/YRESkBlMqY
udoazAOIsvXw1b0UmGB6U8CGjaa978yMcnkbcve4qtpl+ExMj7hAsPAPpL7ROVvv
Spod46ODp674rZBu95FSb5Zm/sWxQOP+HQkzo7Ocj/n+lwdgz4svk+IxYEl/s44r
0b7w7A+pcHq+/JYGH5dsaLEBxOK02rjN3zNxY2UvL4TP+W/PKGDw2mhZYHC2wUfj
zC4FD1/SurdW0jFU0goZ8tavXIaTXDqLqdl9ekvIiCbV3ox1hDd9hQLIJ0YWmkHU
d6am5suOiEN3Sf4bJIFWNuJbccbwvwQGpsX6aKdV86DmzESVM9nmHLAQEEKImFCx
0K7rXN3mnWPaIPCbBK2ObwYBncHEo51ieaPbyB66QlFmdS6lFb76zfi79xjOgZWt
+jLEEDjSa5XqdrwJE+XlvQwLc93q/65hKm2NRNrBvTQlebikcKAyO5AQqHM/o2z1
MFlQaBisj/f6HBvoWCcc1FbpNncINfLrSEr3/wFUAUNxekiOBU3skiseaq+m2nx7
RtYErf+l/Sp//0eBipTZrpsPgH7VwqkZltFfbayCrptsw/GOTJTo0wTc5AMDPCS/
UP+wxDXiYqAZjl6jrGKpOLFo4c728FxSz9lFUBF33XUn5SC4jSPAhYIbh2NmXX0N
KX+Vo0NW6M5AuVvCAR16o5F6VLbrn+SgsQQsQ+y7v86ukb+m8akCu6I8Rt+b1K/F
TYPeriDEDDcVZZJCw6r/mQhXk+tg5agOhJ9Km79kSjKKB9+HIbf4DPBWrxtQtvqr
brsmXhSSmIpA84r/Q39JKBpOfB7TtDqUyN7iXAWfT/j/CPYihM82ZazL7mzPCK1x
6S4pd6cHkdNR+LTBUnP7z80rPdptyIOl8Pw39e1ozbhM6rFVVggxqAtGpFHPYpj3
3MLmBeFOq3secr+kjH4Qt79jatoDnveH4/7pB+fm/qFw3IcwdTOTsSLUb+IMMQk1
nCqboktgOv3KbFMYsqcjWHVLgNThBH4kqRaTpawJijqPDkTHhgfoU83ljkkyFJQg
JsOc8JkTyxuLdWL8LnKfmBAiowiUahA9nWuBJeaIrADwhYfi1tq8O/q26zOMzNwW
QFJBqBBYRK+7RENjOqAk6q8MAOTmohkpEgnNTA7xxK2Zi5YKpIyeBp7U07+0ARC4
YPgNgrIaA73hHmlJQql8aQ9UkJFqXQb5mRSQgDIYTSz410ZnCxJqxhp7v1JpRnrq
tJ0U2FG0ZPaZlpGQrvZ92NxHNQqa7qBneyJy8X/El/ZYOBbqJ9iUrkPKkfucRMdV
Ud/XrM8vfzQIPrDl4n7sROzT04oDck4zw+IGYE8i9/oFJ84JuLjatKl+xuufk+kr
ljgMJd550QTbPm8S8XnCv14tg/uVwFeBpYaeJQe9GKeBf6MZUqUybDshRMPG43fb
ZDdCD282cyzbWY6YDKTPu1zTo3BcjIQkRGYLNsYdxJfdyRhbvRp9hg9swUIwpyhL
b0H5YiizJ1RE2gqnSrSOTKQB/US5OIM+h57hKoAM3JgtgGK5ErqinrFeqfZWk/pu
4ZY90NX4jbCrVUiSW8OjMr9P51ycyHcJlkau4V/K7LASzXICAW6qaufdtOsJErdv
fr9hTjzt7QwCb6cgkvBcst2Zk+AH0XHrmzClO35TlkxTszblDIs63PL/PGg80wfs
5WwKIWNPuuhEqsuZouZI/pBJgJIdGn2AN23h0ib9oIyiQNpHWr+wNQymnUF75hPi
wjGTcv1AH5Hw1rR9ehNYIaGDW0GJnvZy63MVX6DHJuo4JvbDO6NXoFy+FsRVoNZz
o5hEnhTc22XoE/aZ2DCqCNwIm5rpiG4mPpUePRQJoU2ehakA8bPSevYanV5uIjA8
hsXBlsFKJP378uljJWYurBpUk0CXUP6RuagSZLmyRjdXwNiGoIxDwvt2n4FKXYcw
7pEDi3h9XJP9gQUh4OnmNemTRBTi++UKX0LTYMS0iLSlal0clyrtlCqdLc+fQAl2
X+wsYFhN5O9k+CCb7UPD5+7XHJYyCl67sbiBFE83o9QTfGR8NTygZA72UdShY8n7
9bc18KWusPdwCz8gZyKR9+IZzefgQDiuPhORlhVdJu+cRy8hZ90kllD23Ofpbyg7
g6f8dTBxqXCo7fJQZM/SGPn0NUqfPB0yQS/h6e+a3yEbHJY+6OfL8m3eZqo6tpUs
Az1R4Mrm2UQnECAyLJOCmRe5vPqvyLc53puULXvtQSlk8HLbnqQpo9MJLEDQSQjB
Ge7E91de7cTLWSv9JfRLBXqi2D+axpB9BCW1Tath5EBi/3nUvrvTqvDUBvtclTBr
2gOjE+Za4H95t2QZHd45mrIevWUi/K3Se1khvUshN/8qL6r755fNx/98hyiVHhdw
4BXP/QF9J9mdrPXLy5bhVia8ESgiMJ5fEo/GGvbBsAEH/DsAQMnln7vyyjynxetd
5hm4acS6FmCD/Lo1CsuA1I7fSwPkGC7WWrx6H3QJQeU6iegFfAGOksz7aFzWqEOx
STLZ50tLAs6Yq3C5/keJEBqnbHUjrE3QlSJ+yLh/BEhckCbaDxPrTHNZavhSKufw
O34h/lgiBSO1B72MnGO3AGQqv7lR1m0OrUs5gXDUQr3A34VCVhIFalndjQqeBfJi
k86S4cr+BsXqPVwoOukG7vdc+rZicEXHP7RlgLUJp6FycE+igIs4iPQVY9ShpwEY
/6wgViRuW8GK7iX4zm6OhfmrqWUXEo1PClXauXwKF947LQYgI/jZs5Nt/z+9F8V8
`pragma protect end_protected
