// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:38:00 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Kg6WvQLpNIx7eIM//82bMPcl/Cz4uzKPRoevWmZi5Wy7gbHazokxKnXgbvh1+muB
L5XHUebBoimU8EfgETDM6/yInReUtw4fbgYJ/MQsKC/AnLSYSG3NHmbxmwLkarBl
3IWwEfGENIc2awB5NZI6yFXyC/7UrphUnO3BB6ZDX3g=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 30592)
J4dIA4RyEH9lf9d48NZJ3J6OQRY/vrZEvRuSp1KiGH0/Lhoa8XSiVX2MOLi36+l4
Ap6oT6Hn2FLcs79yWig7TijMgARTsVi+1ggfmY7gFxt0tdfgo22p2Vv99E4BLqlj
aCJtIfuZzzuXifVMh0heSpvpunVH93Q8BQc/DLCB9i9ghs0ccjrOFJ0ZkNrZrZV1
XRiYUpqRXjjmOneQ1yFWBx/FCcEoFrtgTXDaHuToPovKAwZsMs/GeZvH9X/F6jMp
ILE3C1A+md1ZDVylOF6BBTSGBVu/EF7uuzRb6PnL4GCNSmuTNYqW+50jfZZ+bvEg
bQmvgeabyLfCm/phG/n7cKQup9bCTiIu4oQtrJWoMTIRxXVFRnuQ71IQs4rVz2/k
EUFGjucl5DWofSztyZXfwsnN56JjUbHkQyelJ4/tgfFdih+TTL56Njk+15UppoRu
EA+IzAPT+lZoS5iBWUGkJgAFq0qufq+QNABir3uyK8+DewaWPV1LOu3emSP3Lm7i
3u24SrrT3tG5bsMtnHis/EZCx2iyIJhx9VpUrBUyB9CU85ijbowENjJlL00ao0g8
N+UWcvuK/1FZhspny4ODPAZV5IGIntnmcFJMghPyNwSzjb0sNUksWQMAImT1YXa8
mdxDA+unl+ovXdK/paozONqk1I7QFNp7WiYVwhbz+cSfpjBHHxFxmrmiB5vU0eWH
HaLVJ52zRAVnvQDOeIAuUe43f/8iYk5BMwiSp8Ry3yiTYnNjdvZ5NbPdxFEvkgWB
GOpszActsT+JRVwlziItQJgu7/ra19FX1q/XrTT2m59qGXd8U2HwrPGreXKIC7hz
aFV9uv6CA1Cg3dFnZZYxU3gWJIvnqZSmNg14qmDLnx2rWayuaFrxQNMKCljq5tC5
4HPYWtOdpMtHvb79FmTuHfBnr1Y00aJ0+/DQsKerHrXZHKJLqex+o5mHsqeIIi1k
Bg3W9zNnDO+rXn4V1f76dX18Y5wA8jK4ALgX/iduZ0q1N5b1YgJRBlOSdiLygSQn
oKw2BVm4Zv4GMHhZ4OB1pe4Ey9V+N2bMpzD78LuHrMTXdS3Wjbk0PJAKt2QmZS94
rKOSi/T9I3Z0aG2kYIHnJZsKS48BFGxyrqpaompXuIdo1BaZ+w58U1C6D2ddCCcT
8sZRvnA83l3LoHEGDt9LJAKCostmCQeCG+k1ChZ6AbuEM+CURzJ5vT+leMe1LtMh
+Za7wtzWKkikv5OgMwk6ErhbuwCDBVWjmOxg59Dt0Dhk455UOjZQyoZTHHYVkAXg
OWHcnCLOwq6sSPg6d+SFj3RC92VM77fUq9lVfrWYTMu2Y5B49Q+4aV4lq0a81Z65
gW5AhnVfIIHV2nJWCb7XaL03ZctRSQRE6nQNxk/4558LdLNYVQi2KSx7WRvWzWT3
IlKWUP33Uj73r+wlHFCkBsKYzyUaEXxNQN3efQgOHNQBEPFm4EeiuercOI8SfQla
QlkdF/5W4C0Glt+ySzv8Z6PTibMrqsiBPaGrlNBBVtgKqkDqxYTBMPpa04kbII2z
IOVkweB9d/ZijK+wbtipCl72mmHKQS0eriDOEkUjeXGZ+qbwQ0W98G3BPBAY5lkq
EEJphMRID5dNEiBxAqRHXCSWa+VXbVN70w2nV7D9SRbr+5BkUVJOrLy/DyCsOUwV
LhNqorhDEh9/0uf9wi85C/gUpHJVns30x2wK2Ijsc9peOo+hcdGNNmOnXas6xKsO
+U1ZtCeqtr7LuBHq2SlYyRwxQn1Dr3ESrnaHQesquXDO3qaiwwJ/54IA5BHcNSXE
XGxz+XnkA5Gq77D9NOAultsBVMSig51QxKozFq8N273ychYAbF1E1O5Ing7JbIJK
+V6aGkXzmYd9X400Q43Blqz4UT0uWnf3il7rFpCjTlzmZj3eo5uihoSlhd41t26Q
SZcv0C5PH1IM9EjiPVq7pRwKLtZyYYWrFlahyR3MRlzimT506te/beupEgGhNCL3
NIStNWNtyfZZl3idaUYrtFqYT43fG0UUNNinkSrQMI/2KrTewCUwogR1cpIT7eUd
iGWnRBLIrbs5zDUburn6jDwcJn2f/cK8G1TLDJ656QG04DZmerxJD8WodMLxX/ge
SQt7xfrQi+VlYquCv7HrCaWW6oyQ5lTuBAd15kdAMn1S5SXwPDc+KCVy3K6cSGIS
/4l2LsNoUM0SkEMiYquMiPxPKckCiVqusDIzWxsJ5pASwQmaQfCLuMoBEJ/pRbR2
FaxyUdblln41cryqA47d/0A5hRvJV1WOfjTJElF7z1SAfLtplXkr8yO4lyQLMVBh
7nBN05DtByniOejOz4lAs4/HTT0zvbYfTmh/tM30mLF7Njpolujhcn7OackpBKF6
nVqOUGysdrt2HimInRyqIbbylMSMmAaq1wIhHJm58/GgPlITfNotUWBi9BrE2qZG
ujUTt7m9EpyqSFwIQpeH53bxvjAV6etsDyzSRJakAFdMqN9+vdtWrd/l4vbCDxZr
qtboJeWoaYYghsQo3HZzLZ6MCQUc+zubuLRFTw8nGm4Le+l2/FE5IAVM+3nUbuwK
7MpLoH3k/GP+A1b+Vf9hU203VoHeQCvif6GcDyMToIN6Tg3ewpTuMsKaB49ySQIf
Z56mKBZokd0RGaM//fCCImrzQfw2M04GtCSz2LGy9xb9bKBiJs12zvnWFQkQc4ld
LAHvjgAF5YSyb/F5ODvl7ri9cFqz3nOY1h5bItZqAwaJXHiEmZ9DtmTpzDXMOtJY
bq6GXVWo+pJuv+/Ilo9u0aE9nwDqGUMe5xiWcaXKAzW4Bx3vg/RB+SeGZw4FZKBF
HfsoKDUvK3vp/GJFVXs5cuq1e1p8skEmmmE3x+7tJDrMY965HHtr60qCv2QE0ufk
d+kKS9gZ8YqcC/T43WZseqHmQBKilAjtqFj00f8I6Nf5T2YgcRbnvzs+zL31ieFc
oNZWueQYoUOJ34Cj7KHZj6tFO3ydIUej1+PPZnhQSu8ORYPG4EfU6H0JmoyQ4H0L
Q18CtQFfFd+w0hb5FD1MsNGEuWqm9IeWIliIf22f/A5oGBMXdcKqWqwYo55CIEfg
MuF68GcOWnoVOVaHmEXzlZn19On5K4XA1mMCVZK4T/R3l/LdZyxWvKF7UrUUQx8L
Cv5xwI3ikjw7HKMidlEKVrK0e0X3xdnvm6PE6V6MpsvxN2beZ42LYeigBY1IszsG
qyKOia1cEoUMXazZBU3L3LLCiW0G7Vi1DBel8dq/yyrSf5K3mVCPy4t5uy2INSY/
TdwcQaoC318nS5tTby+0ob4S3HHhjOtUSI/bvJUOfWLaOI5+OdKB5c4UNIlDIRQS
x+rbUliJq2oRW9zy4suLTCy7tmDO4uyke/WaHm0H8Qq3o+NspvDPpiTAo5m4pucd
CT0erXhF+Xtxkegixx5oVA1Ys4OtQlMvQjA4y9tPLV/1HjJqVWztySDvnK+diyjS
HPVfvn87OoYTtXVhMwdzPrJUaAu99d8/nodBYfutWNYhliaUO2RTtTB5BwfM/XqX
nXaVo0cESaiV817A78qy5xsRf0ReasoeV3ilPvUEjYY6qHuCqII2NLwjKsx8Q/yO
A6km72F7+hZdvKsGvm0wBeNzC1zpOTy3bQnOg25BNVdEePSe5mf7nsgLEsCT97c3
nL1N6cDZZoL8kr1iXBEKp9Q2YJMDDegRlIWtCDE24aoaUIBbTClQoCDi9Jdf3Odm
aR8GLdGmVhqvpLgpTpIM5bIM/d7LDJ1NEuXCswg6H8CSGY+UHbdywXQ6gTFf2Ha9
8az8KBj/wlJGIZFyFng79REXoSif45kO3w2nJl63m6zpIi40nPmAdM0qixL7Ee3t
FtkUwYFxQse2JyURFUJ74JBSNQy4UiDBw1xSlROn6Ef0SjdH+fzS3XL0N/s1Lj3V
j2CshqVvLeYsNV/cpB2wy4c/4flY6nwsWSbt+9HsCpn39IRoipzU7CKXBZFU8sSR
bubg5ENT46ObmUM6umEU5iDJV6Mj+uW/EE5YV1T8xXY4ZfSPYtzIQOxD7Ec0T11n
qSSfaW56/+LSwffEAgJlmR61N7GyOcJIzMQ8eYsbGuaGZohY4HgTVbJPRRKzQKEQ
3n83yQzUPzsMsUYPejVmrgzpk576clAOgk+ivkWbgSk+cRx4qTkS2O7RpAvk45M6
5DJmBWUf4Iu/nUV0ZvnR7HSmUddX/oAsPolm7qHxd3Bg11gWr4oAg6XTEYoDcguP
tpoZgb3emk6GMBVFwfc787Zh9h4trIHYHJZdD8JE+Y0os79H01U8d2W0F4nLT465
xlicM4QKOPPpz7GOHlhTaO06qxmXTgSVipvHVweFPgSqbm5MPU2DtDDjDv8tUJBT
9t5DvdNyVvyhrEXgz2nvnJoPQo2U0xzcVzyN2kXWhGpLo8g4WR/I0EnLPl101d2h
zCpg5JzEUt7hyXDgpWWenKsGe52KXlabzkMVHIirDQluYBJVEWiCZ/DwilMqTdYv
3UfnoTZ54SV5LdKtphD4GrUSTuhDIvbVhn5PaIghyaYnL+2naPczzhdmfLCwZVPR
6M5oFpqrXmq6mEM1QYFE3l9fI3dmiXXzuX90YF2Lp6WDJFcPphpdBnNwv4KZ9qQ1
dH22UMlhpIwGvngcZNNkrPIv45CPl8TN9Vlb5OuNrUsVH6+DGc957eDDTFAR6mq7
WW2mDjsyz6QEzpG65xNpT212HRfVyYQcUNW2YBNmI4QyhHJtQq1tLHuN8i4vDmYf
l8O1NaxR2RUbUZ9lJJloFybto8vge6rtMuRV71nAvb/JfUqy8fbFuE3N7hXpIUk8
jKD5XEFunJ4fd1h5voaIcx3E2ib9/6hvruuhgzqjCtngYnRorCC5BVaZd74/52k5
o5TYrXo6B5w30UTPbYWiMaAadHiQI4jskVioh8uhLT8th3L2/L0JW8S3g1TB1wes
yZLwyHGX79yDFo1z9ZEqwvZXo9H68tq9+vZDIMOA8Z2RPsYxqPzbcMVHqTF1KUJc
oIyFti1ZPdhNXHUnK7saoJt+9R2tlsW8MhFZbBu1DvZHx+FIYYRl9+2zGe9RGOSG
KI9NV5b2FeKNnADMXOKX0Wu35eb0RI4xenEeuLh7opT9guIABPCxnjACxD4OHfgA
CVK17hrDMb8vvyDktm6XYL1iJMAFD+HN/y27YBgK16F+bdXL/9EofsS+TmpCByI2
VmSRGSyQUo3kRGEHuTd6MlqQO5gtHHVYS2o60QGNsxb13aqpXz/uyg5k0Gg/8WgU
xDdtvRuGSiZYBKZD4RNv7Gdyg6ZEs6FZ6aR8Efs/+H5Dg9S5q1jbLqsaprreTY+x
kCpeL9xwthjjmdjGXYnI85Xz2HVa+rRKPvJ2XERkE+md2zzr0eFaQFfu8XwgbO30
8jVLQTK6u6DdPySZ+PM2QQhlfA7YQCwifwg8yCXIGncxoAfx5ilAo0AVZe6gi8ma
At15ey1LF6KmVjMAq5Y+DA9FFPyAZpQ2MssZQ/hcMuH2qgNOZYeF6tPATaR56v+Q
3FZXM7U6CCbAcXwEbXKBGI6aD8fBzXMeG0OWnAhj5SyU5v5ucyzYZgFrF2JCt8zb
yi1mub/m8QpORfqcVJJ8vGTaXlvRt2cHfdkxJhuiL/W29c3+wJlu+uSZezuHnF1J
TH5fk78agP1DLbh9IZTVsRzErKw/OpVi076GgP9ZqWjSk6Gn9MoRoa4na0kHzMUt
+N1q1ryzkVDWW+bYpeMd715gupKCTC9y4sBS9mc+uagrLNYtSfMqIRq6Fj5eGgZw
OBZeY6z3l/3iLIwMTI6UfGf9UKRbk22iRVLFJOFEnxHlTNMlfi03KpHb2G3qA4sO
LUAfXZCziHp5NAOQrjBRPe9Do8iYvfUVlCqSRVKKymaBn+bFAnQ64MMwglUATmbY
cDkd9efR1xQCuQkd9ete8a6jU/TE8Irlf7sOn2M/2p5V3hDGtw99JfJ8N/Y2JokY
CuNQQgon14lFUpkAarM5aj1qcz5scE1q76sbBvXpM0YlNbKfdbUwyw3CmhLbW8CC
fOc2Tn8lylKfx0OyopUr/D8iJk2jrRG0/v6yM1PGCshlvnFfaYtDE5IDfzNgjz6C
MhLsHeVCLUFlyyCSkgYBuASRzI7gtvBcXcdOgUFxo/KOPc6qiuI+lv83DyCOcDWv
q/AKtFvOQi5RF0o8fxckmp1KUTEokVlRWnOasBtxAhUFdEUnQsqixKYEJ7+BWCXR
cqOD45PJy2/eCgIHspJuDjZqdfO737NaJiOEjpvbMpljY7VvNKitU64MepkxeT20
x4W1pSXfvQ1z98nQv7V3JZ8S7FKDMc0hV7h6v97Iy/ttRW9XlOtesq4mUNOAzmFk
VQcmJTsnMhOgv4aQmDzxIRLE7m7heLfPCbEW2gxGsq8jGG7rVz9Ti5tPDqxBefwt
q+e0CjFjrRio1K6hoRUiXyQYf11vsaiqrlFoO68uF/aqLmI/KpuMdZJ7/NgFofYa
vZiS6X3BJaxETz3mVibfgF/lqAy2Idi1PFNlawizg63Jrk5dyaQpqczH+v/3KemV
GdTpLA+e8tvZvlK1inXU3P3Xcp6E8UbFD/q1Vh787SVIxHsKTJJEc+Mqq5Zw4hzn
jl3ZtdsRMFaDqtHj0lrQ8T5QDY+qxOWjjMpQ9VqO3PeQYulZ4ZoXvRdgAzvEkdOr
Kb66lNy6+lIBme0SR2lV669U0hKne1Ip3/7q/Ts8KTUgVVlWVu3s5YuQ13VV9icC
PnDN0EIxqEV+Vu/Ob7bEiYfb8qhPUKLNsQpQKtr+qAPofH33+w2VyhJG4zVVmAib
XFF203BSl8nMzZEXVme84ASMOwuxJU52ubXIfrXNnw5LBkD0Kqpn60928brxKRSD
5uMgHH6bVszn+eDkkGSVjEG1IHhfyK7b+T8F2X3RPjsRp6qL4M+E4TkFlZsLaW+H
cIp4Um5kmMP/SqwMHhOVUuJ7nxMoONH9dQCejZi4ygxqkm8gaa4csA0pVt7mpMMz
AM2r8tMdeg1thEMSR+6FPDB8j5G6XWtLE4eyPAo+FRe9k3njmvLjPeCfZrtTVAn2
KDyg05UW7azCpTqaEDiDj1IFehVi7B5hCdH5hrE9+vK0htt7qLXGXhUUW/1l2T/u
JUYKWdbaB83RoUKhKi74UOXOUYHapRV6TL9hYwpaVq2aktHXNm3FSnoliUVzNuJj
CZACPOFtTu2/lCES+AV2xVAQK7KILPU7it8scuw1mJgKzxgzH/1Unzp2gAPbhpZZ
/ZrehyKfbLKuT66pVc8FYsCoIUBlREey5UzfntaUyDNQoB8R+JzkPo9FI0KhI4Vu
RIHYhZXTkIQIJbBo1M77hZ6DjBjzzoXgnN9kp1xz2d5nMGHQY7fLTJuUayp7la06
zZoNt7AGTCRZMh5i1QbsHefdbCWdi2NjdZb/l4aiOAeFPTzHIgRHRI/q1GIyOlLi
HbvlSf/FMwL3aIIKKb0nZ1CpQAYOtaJ2TTCn90BPBCLCcpj/9fvG1w0yU3OtIKFo
Q52o9YA2YoFzxJb4thkyMtOnMmrvpNAgL45FUN4wwChWKQspHrywhW5J1+nXEeql
YZvH4nJlPU8KDqkLlMUhj9cjO79e7Boig8NCvCd2l/HTTFD7gakqRZH/Wbl1dLW1
8YT6sgQFwiMa/ogAJhoPhmH3ed7qZXb3bqzQFDKGRbhtfS8zXoYDXd/1ap5sk1Yv
WBpnuVUoo9feWSkW75esFdiZb+jqMgN5P5k7diUbOUoKTMsVzxbEjq9q69yIhB4c
iIjpGDnta15zVq1u9bWGC/dOfr+jtaB7fe8Cn3/GBcUtIcW2vsUCl6yrfxCAsCXT
HBH605CIoHRuNTxxqOmKloB9RBcTJG24n+v4P8OoakWow0QZAsLT8Wr9VSuKGUz8
75wLH1hEiJlCOpEBlE49yFSVba8oVP0xyWIdbbbm2MSVJCubdv2M7t2Y2Z3hVyVv
dB3xYXpjCABFhjrMinD3m0zcD1Aro5/qI138+HednG3WXVziAPQFurkt57CeTsAQ
Qzp29+F8j5zV4JMCucuMjC/WaQjhU/Q6M3wesEwqc6VBLfbkeTlTT9tAuGltyP+5
ZE3Cu6TFLFGrBUYOcAJNVIdt3Viqd4JA/gZAW/cQrNJERbH8fftCLsthexJC86Mv
d2mDdkCfp225YnBXAOoyL/xTQirLfXe4FYkEBKKfwHIYEFYoiG8qpFe0hlteguNd
b9tVdU4SZJLNHbKGRBBs21CT8oAFbsdEFMyB1a+5J+Toz143+3X+nfx+9PWOR1Pr
mH2rl4f+xGOgiBiLUVarZU/fXV92PR288qyPiwjwCLw65a+AyMk0oV2FkcWp4gq+
SV7DSK+wByAdSdv3qQtFXJhJCgNsFVj6Bgen6KxLevKaPakoCMDKsXXPNrncchxj
lHo3jCkt0VzJLnfZIJlzrA93RTEUM7mmcYJ3MWzTWAmqwZsGCF0oL8wlJi2MyIZk
5xiaBEbP0KzkDja5xBFNHd7e0AXfOVCaa9IVHquQ+mLwKEjbnUERawZ7fl9BQi3R
yIM9Cyl3uf48ltMBnaMd6PNjxbZ/PxmhKjFDaVul4X5agqWxYg6msBNMQQ0jY8lU
wUUxEQUOzo0V2NBV0NpETm+XhwFvcMnepkFAU0btY0BaWfGvWqGSR5MgWyJAJv81
bSQV6NIhPldpdh1eNntTCc/NoVplWDl8Vn4/0XSFo+2i9FaLkRK16Ue1XYn/wXit
0xb1syx5q2MpJj8RO5MZrH/dJTQ3gSI5JfieiBXuwLEujlw8Hl7VfGbPhssmwYs0
qdK5B409e1z2cYG2Yi9MJC2ph0Pa4d0cIeKLP27ME5s0QYOYSYKdO0RmHZEBrAW7
9TGR3pWdu2EbL6sPxyv2r9Ll/k5NkJeU1ptMgTp8JsKfqO5eOwcGZeug+chFJYlZ
Xm/eowUBwSgv7uXTyGC69Svt+j40tIRZlQHf0iDmchF37vP0RQNjnQHoC2BwwNb0
XW+osmEGT3t6VFYilA+8vpJR4ED6yUCPThTOj5s28mCBZWSEFzezOXI1uNaqUrTQ
JXDf8AjPghmotsIIu+5tY0Gs5pkTJTDRFALhZMprRSR9J08QUNQHx3vKWv6nNg3e
h4V21eGv4M5eaNbxDZr+cxwH7TdvE1ozq3kLwaZg+uFHiLcaJIiG3WjYPsm6sbxg
RpxAh/uL5LkpIw2QNdRtMJP7JNcNvmTXEWnJzBLlq+lAJac+VhcZWr0efSEtSHoc
DkfO+LHt2U7pPGFCnDrqQk5evwlURRdmmJtrJfEnPpqBrXS+zIpeEo+5kKClCiN/
G9x2Itkki755dYabJME2jms+NnP7Nu6xhWwnqxQQNGKaqkm3GjQ3fY4XgMVCg68r
qinuVmo3Y/neJPZVdg0cyR+47/hFAno0u76/7EUV+T6obvzZMT3ELSXC5kKTXjEq
CHgd+Ql0r9+9+GfeIg5ClPJxZ1tl6+w+VUVKXIIrq14HlbaTx+Emkv0HkhX54Wt0
3dfGroPygs8ntt9+Dm9qeV2wlGj/3J1+LzVrcd2kCk4ymS8+dT11m7ySQY8QkBZ1
h3IKN2lt7znrU24Uq8SELChp28kjqqI5PnFMb61qOpma1YaWTMNh0OnUhbAy6Zt5
MQPD5+ZdRHI3ddjVNGAjudLVveDl3+D7Nr/1cuMX7JHzyvWhLaymcafZTltcH1ps
wvQfOVWNecGjQNvZ7s1VBZhAnQHQG+2cllHvKVhEWTV2toVYpRwAGQ6GYBfTLzxe
A0gNrIL6cLjLduaF+rbeo+rZ+kTfaar6oVdgrVsRUfwnS7JtsMYFFQDPB1AggIN3
BjNCtrqcLyuJ31DbygnjoJG1TWSvozyK2+DCPfGMohY1l6wX+4YkNoOdQpaZjslt
CQZC9D3qbypRxjD9WnB3p1kwASVLvd9MZDdPw5iYmQ9hJpSfF2cDUoMEdITtl+FB
Ipi72Ddtwclu6XxyvKEKgS/Uo7VSj3v56pKMOm6YDJ6Cf7QY9Vgpj2cpS87fjqhJ
izlBdZWmfxv6dDNWUuEeYFP8kA/BBQ056/mzth1IRqBbNWEo6MyUJO/ZI+WGsFuk
cVy6au3D3tpcjFUlVaV+cx/jWEqgx9trALqh8xu0KrinSRAbGDrnmH2ArlCrcoBR
3/P255vgdMBOZF5ovuBhYeHEfgQnW1e+vRgTtqlDT2ShnNOubVAqLIRgEqbnT3VH
N/p2zKqxmeqdWzVdlysMKmAbe+2q0ea778k22NS+J3cmFVyAWLjb7H4UQgV59ri2
CWPs7H4gydCtDD4Hjzuwb4I9wDD8W7DlHWadH5GC6535ujkXzWahyxW+oCx0gcCj
EL25XpHNkhtZGmxskQY2LatABsO6Kg0pHRElBh8uCXZFW7Qxk4bLvMIzqp6JlEOG
H6zWEu+RSHRQJISMeydM3RgICUzG+vbx9Gz4LwV3eMlgRw/LuBtnEnjfkF6R2RO+
OjTw5pEg684iAELhHvT+YBr3KTDNr0Q8BlNqs8mgrd2EsC2yfQHuyl/6rZCpGaDg
iRHbS7bSbDbu9M9KHJSqfHHXRnQViMwIsNY/hrXOem9S0+ama5TO6gPvp+3vdnXc
pz9zcCyAhxc3lZnXWc9E93X1gRu6imswUonmUBBnklNjvDaNMV5xA6zjgHkjpnUI
sql20UBWsCA/cQWscBtSDzk/OTfvMBkREfxA5mRhm3O7P2TtJYMDAwp6cLp6aZf8
FFq+e6V7yOTzToUD6ePDQ6K1lFUEoOnnpl8uUyynVDIb6nUJ5D+NqXa/swIx2bxf
HoBBkVZS35MUHj0FfgxuTFqNL11drLAIITmuoykPoFNypMdasJkBaD5enPQqfRpS
GTRk/lsyeOjRL7JK+u06hznzdNaSXCdXQTsTTNkVX6ajbEejYu8s3LXcYoACJ48u
dJsE/XLWs2guhDIDaCh/tzsuvWqRMFfnvWhaWo7VhRoHH1mYGFQP8tCIqAZYkMW+
7PABuGi48AB4urX/WoBYRbetyKfTUw3gbnISGVchTQPgtnqD6cmm8o31PVIize1T
BDSqiS0rJMEQX7xCuMsShRlFsdDYApmNqwsfvZO0FfkZJOhqf9cjop5/pAtDcDX1
slx5twYfimbeq/giZfTq2wBCb0kRBN8qC5OlEHSGYX73o/LHg3xzQw9LkbkUH3/i
SrEcMFaqf1ZjRDoRQtGtveyIRZ0Fql+LZb7jpHVdaT4eVKKBD9APCuYS/pHkVhN3
aMuWiGoLM8sbHO/gxYh+zHh1F8dsCdQ1vMCWWuKNYELcSxVD3xsA3XH41omE1n5G
WW4fKDhe76xFw1sRQ6gWixMYTM/BSxa4OWcPpEoaoyBm8hrUWCJdXZEYF4FO21Dm
SOy36A2acakA6OUYOiIl5p/+EeV5R9Uk0ZQ5nBtDpORL1SlsNtd7GKoMbusrbDSe
WbHNrgFSmNLsR3BuNDA26cG6MAV2B0ScvdkiGNHhdQkxo8opg5msEV0SQNKdN3Tq
UR6HgA4AU7h1lKDZoAsjCoxocMNQ5NC77Qw4++SHOZIyINw07wqrOdw+tVmHIYrD
ZfPq8c94ilrpSSfSbiLPZwN2qrqkiu8rApj56bs8daiW+Vp8jQiu80puzmM1jdSW
t4zOrSutAZ8P8TRvBg47NMmicKqWeknEATcpz3duYEatw5It+BpPbembw603eGWz
gM7eFUdAz5HRiFLaHPFNsB8o4ItXn8SP9U5jJTuJVCnjDjQxO5GSRb12dI7WKHUL
4U0c7AePUyJU0HQPs4aeYzRf+KCG+bUMowyqjjtecqK3icH6GMY2Ee9KPYFH4dsM
RQ5ZJCvmOHnAGMG2f7UjyRT6trGWy5nZ9KdbT+ujz+zD81k4QQZKJWafhj9ljT6l
U4CAp5oqnea9ywrdnt+qHUy0oDb6d0VJCv8sadAsyrgZiE+QW+aQI0T0PxRw6ojL
FmyGwq35bjuerj9O3QPpPvv2W8TaxDEOiHQVsQPEiYuY1Sapoj7Z8EncOKqiIn2Y
EngAfvZ2dfGh+NlgyE8q3rmFh02hx34z2pmm7LZA40zfxjcvKcgH7q6BuVCNwuK8
po1J49J6RqmrZZl4F+oyOv7gvazQGbUDN4I9TygMos9HLTjyeVRDInfU+f/XK2UX
r3gyx1oKPvueWe1k6PkAp6PrsiiT74qbHzPSITm+ABxFHBPA8oKFL8Ixpr6Qzpq1
24pSLUvvc+N93hZmouO1CmZLE/+2cWofrzizRFRlHeT57q6MpFWwc9ONoz9Ckn0u
LiDiiGvOs35Y125bAtqZvILjPBkRfNuDIz8yQ6QAHpFYz2fAdm5M5KztLO4DU8Cz
fUqgOY2Mf5UqnHmAWjgzYP0lMyLKkN07dF6aRWVRV97yB+zwk/iS0TGlPQF2yNcw
5BlgQ46qwbjNStEro7LLraBt0KLZ9OxRdINU7N2FAkB44p2elVLTrO0gh7nMfWh4
fI3UJGRuuNQ1t9qbFQnu7XkW7gNpCgeGyY0FdMw7NBN3uw/JOtsDSGpRXwf8gkWd
xMwp8F3h/Nxsa29VWucDwekz9CQvDMtxWn/6ay5YrATrFlVc+5k8a/CtGbbNTM9g
diGf8rUoVZz+fPf0CO/SEA+sZS2CPea2RdbQbAGRDQVbACPeKH1O9U7M1rULAoDo
qGMrfSmkahs6FBXNvysAAbItGIRXn56iWQ1Bm20YKkit1cji3XNgC4swODVHcbHl
LL8q0HSlD8Upngyd25QW41738+Sp/LtCBBu5xCp5cnzMfwgnKU0kjNOXpxUINOwC
EUeh63J46gGRrj1vCuBuXT2n5IsSz6lsoDUpUxZM5bJjM+JoFNl3ENzgwTBEYOrK
lZu7QNQkq7b0+PXxt18+oI+W4JxkXE1qcg1oOTz+8d9bMyOO0c73K9LdzPKXWdwr
T92w1IX9C0MhDAPL7nw+SN7b9AsqFhX8OhcCAL3jBojz9DeH85xaoa0QBBEXGCq1
DvUXdc5B7+HxLrDBIRe0MDF4gZ4iky7RXmHWtvobe4rV9LKTL2C552583KKyABrG
EMAuYi5Gb6qT8ctUk1FcUWXjq33+GCEm35LYlRWUSsCZmu4VEo8gy7+RP3s6+vcb
eiGXwbmQv/z+SW+EH5RObCNDaBS7kpiMgYtZMKoUe+3JLBDRpW0eU+UaqHPd1gFp
qbs5x4EXm0CrvZfk1eMxPYj6hvSEtfR3vq8YypX4ZhNMVb+REgaxO92gVxDHIQda
BE3VZc8GPb/KUf4Sfm/m7snOuw0hCPm9j1POXqnPm89OOyNudLfI4zDVqZXWRh47
+o8GQQbpM/D7aGN/fqCSnhhOfnPbGHobIZcBKFEuZSjFOP/gOXHFyyV+I2WQpP+J
U95fKOs87M6cDNIzy6RJtZs0top6dvEfF055XEn+E5ue97GfhJJwyVhiZ7UV0khz
xHtGbsanC+uMcgzl0ULl2bZl5+2TIgPx+dg/4DJP4LW7lHn63H+KiGfBZDaixlju
KfWAJ6A+grYSw7lSkgw48IS/wzRXOWSGRYf7BaWHeLqQIKFOYlb9fc/h1JUyD46d
isKFbbHw6mVfO4HN9m1CM+ku5RlITnJ927aWl5rfV5lJodpfMgpCWiQwXidkXe27
3rEXGCG4+dJHQsj8mSTUVA4RtTkGph/tCUGVqArBeq992Kqn/vs6q5/9nLmgA4aJ
pXhfZINNJwvzUh5yjDWO2MOfQrX5YK3gQe8GV8JvatqTa8Hysgtlo52VY6bVN9HU
OM5qWgWzAIdaExY+osUOGafZDw6j+gdTeVxQQUlwpElfAicDsNrmBSosg0ZzJLOy
NTUUJLASGtdv+CY0eBBAwX6rPx4t4x6do32LGNBfD2Z98jQvPvMLk+/B2+U28Na1
sfVUEZJQNju2JxARUho/pq2kuuefA1kOVwaeoVSk0meSYguipXmkV9ML6HetMotU
kU2IuKASqBD6yFwaCezACq0mCKnkTaE12/Ua51DjeqoBMmTpwmEkXrlm4+vuLfcM
RE7+bjWUus6bXC4HUqk7nPKgjdAKGLJPmyHwQZFBBX5yQz3D0XExkfi+/VTb21cZ
re0Tvss9aRd9QnLaaB7nKBkREONNoOsxvhTdnT7xeH3qowzvaRxxc9CUrdEhKMqV
t1eBYfWdoblVaYjqEYtGxaEVOpIqCZbiCoBx6x/u6CZdDxHN2WmuSgHik3TxTpBm
SVzI12E/sZvKPf2cleDvzED6m7QBIpReSPrVjcGykMJDCPs9Hclj1j0WWABDRuwY
Hs1geXzJdozJUmjw3pWzlk5gw1PdKxsfxQj9O7xFxUfYEASHFAuf39fFkPP2Lh1l
mDq48sgRQxGweKvq/T54m9dwWzr/xNQjUpYnBfjJ36g8v0QzMAfgte9nkUGTwy2r
7FjEi5GUdw69sbATxveA2dLi9Yo31DMfY+gdyRV1y92Jiwo9p36CGSyN2KTXmFMz
ddcmYbPAr8eTmOCJRDu6l8VWUfPJzDW/526lxVEk75w/ghc785bx8CzacDi4fsf5
CdR/+lM2Fh+Xr/4GQoXqDH3NEsMT5yawTMGJ4FrZkFIGqZzUemO3Hz2awB3vjxqv
LbP3f1RvfqO9xMLfMZb3oXKhbfWtSoghmre2Ae1OI2IUmtlGu7IUJ9TLQ7sKMAhm
JSNB24/y01aXqX9QLAp4yBIkACQigAZUx4w8RGaR7IfeCed0Mbfd5oO+vpR7C9Xh
1lvWJFpE7ZZ6wOBU/ZF0c7AcwfZwodYmzDfdXLTQ4Vk7NuHsXhdxY4Nssojxiqnj
/uLlduS0SgsXZmDl33VBsZitYIcnpyDo05zjtWcwa+qqYJOGr6PliGpfmpuc6TuN
/AAVcnmXJqTyZKcngaBJm2G8wHo0mdtPxJMg/Quv7z+Odbc8oxsHfeA3foYPQKsm
G2/qR5YyIxBQEHR/WTUAjWxutIwNPGZ5C8lNCBo9+aAqkra/ExsbG468CWdgS3o+
NROQgW5xlb7LhomgV/7CqdiD5LWNu47Ee571k6LpMsO5f1LLQay0+yM2oluNiygK
ZXeyuzdvci3kjKSjci9AEe+Nzsry5YSriz842axjhSm7ne/r9Nn+CAfO2NkrcJdE
LMitzdXsEVEYSv+e7+liL96O/48nv0bgXxWx5jt288snihIZxHn2ZQFjr0zNZWCp
ycGgusDcS7ZPLwIj4Me+L9C8+hXv6sl3RrUoBJXd/0h5fu5UI84pZjUZvftcLGQ2
ZipCQdVEAYcSyDd7pndgdyXvEorjvq3VEePoUuwhoqpiFduvbsSMGL0gXc0SSSQq
l2d1sDKp5ZsRMnzGxvJmhsO7y2my8YTdbpwBaypHdaoWCTYL8wLuMLlps4yrFf1w
jkYQ0py+8qu/pr6ngSPyXYqGgh0XztgUIPK5x5qieOz9qTfKXOmtLebksLAwdQZI
QI8uKPZt0XmrvEX3ZwlPc62efECpmjWG9o+pjvp8Fji27oMZRWDiyCXR2NvCI4X3
y0Ya0Vvnel4SpvTZBl3ChI1c62fFXmeeC08ZCzHu9SXqpJiJyBj1BTwEmYzv8TeR
/InWih6zlsjJDqNiRQ/8MGyiG8+h++U1VHtdUkZgJX98BcyP7bNZtzzw/aLHs9J8
URKHmwuDCViiFTVtx/CBfDfBSsqVJdics453zIpnZWvPl4d0gJ/vyQw6dpBp7Tms
YSNaqINg+5xP0VDWMb6J5dFKV0OGRs6HTUa/VEh3BTnNns311mcICB23QfBoMj4Q
Jua7blnbPgN5dDH2GuezwUgKXXkMZbyAIDlmbnmCgWYiv6w+1hgezLSPsFVgfUYM
zxWQLP9VIO8Z776YVn/rX1PowzwL0V5nhRgaIwBw/Ix495eLGl9ayN6dsie1Ipsn
lY4ZDv2AjGHkxYgIXjZma7bl5Q+iGUu1HbxcLYRj8j1dPrJBZs5IT3kgGoWHVV50
NsHR+lCq5hf8jPwNqEDRdRU8qJ+OQfDDhHSwlRTEB94OI0rbMqbzDPPX+1LiEJCm
LmHJdX4+R40RHCBUICC1lQKiyIFHFfqQ8MVnw50A/w4+XTQ0SDxGo10HIntReRuX
jkyTN/u+mPxvNSUVLjqioKFhsdZtLhC6JAmwecyb2ufaLEKl6TR++HAP7n6jvziX
x4BCD7D1tmabJitSxT+iedw5Gokefq2fhoOg7UmS3nZFtFI6oYvwqQb7C9ipvzW2
0+mefonnPWicJanyw0taHs+wdN1JaQfFEY5wTt/ZbbktdDFfwUqF/tGXR8aNieH/
Fy02nwpqKIqShTIUR0XbWh/A66/CaE3gOYjr5JiCLhfF2XM1XXSpHjA1XsEhWB5f
GaJkjDRzIHezXrHq2GVYzz7AembYbqHTqrUL7085Yy2ETW1qq7NCIjJcumOQ6jsp
021NQ2sFgveXjlFMbeVxKWkpPAT9IgF3cQjWaLNlY4yTS8U96rwbWD1oH7OkvSEb
d+2fPppOlnQsx77CiEz2XPeP1hn7YeVBmFGJKSK+58AV30TfsC/VI5fvX4aHrjop
I5HnO7aQQr0eXWpLoiqBQkFWzXNAMiYJPt3sBNNGMy17CrvyOPLKjzoIRjCCNXeF
Z/DE+W9wBFcD5ftIVj/IzNoZwF+8nzXe8oEeiKl4xjqRaUSMIj6TvTPf8IcBKlqI
1JAWhCqrr409fMlfbkw1aEhHQLjkMqMJsbX328HEBQrW0A2hMS/Kodwsfku1vwgj
B6k3NxfMLa4FJn/8PFelef0yjR0ktwTPlvrjMQ3nCiU9JRg7BUq4+0O3L8ofeIRB
OFkkiQBGD+MzPwdRW1gbB8Vt9Oq51lqnOxtWaguoSt9X3oSUpnQi7bQMSGe+O3oC
5CuuAQuo/a7VpM5YRxAoMW9uopOz3cN+fraS81pL1rzQnzSLxTb8eCKxBeiShOc8
egolmAQeAu9W6esXAEHsbkzc4bR/GAKSagmHyRdxw2U580WB5iB8AYtWiMcLHaLe
6R3Wui/CVesHvjeU/0NwBQFEewfnRi3cubeBO52typEadiSYH1Oo76ZA9cBK7q5d
odhbRRIKdsiEDj44h+0oTZwPSKS1KamOShFdNczzOg5DVih58EuL4zMJNvl6nVBN
4KHTPszX4OCJ9cNiqhj/V+B0cvkfyXHDPSmpFwlVBJCYUcZhPbo7/F8uqB0XWNx4
0J6A3tXgnGARm8aTQNLEKWyIvvlVUmZrl37+CmGUjbke2EgfBWusEjRVjlSqdqR4
hDwR7DbgttNlPhRQrPg0hKginvRtW3IXI4sUsTax/7nmwTLwPJBglXyNFJuB2EQA
zlF/byZqW4cMs8b6fnODo6AsgOs8Ewg8c+PpKhEqAJTBlIPrDwx62qhNCuvco0k8
rcpUhfcMN0FqO+S2DMt4IiD7tJNP8DQ0x+yjjlvy3d4Lh0ciyo0Cxs3NbnpkYdw4
XsylvB8tFeZP+EOk0w3+tKV+W+2Sgry7oy6aVQPZ3EypRVrPqFhXhmy4gZR96lIv
lOU9uxbUwl4ALN/Kopvq7M/4N+h1dQZM6tGfyRswBKQvmPzb/pCHSECPNzkXxx8K
XG1WzteNx6mBG62iDi6VvM3wyz34jKPcXSQoxYmYsEmcn2m2eecPyLU9CWkoftGh
AluyghWHAqtsHXRvLDSJbiJgxa11mWeXbDQrTQ50oKxi2EPxW0/1XHuAU4HPCDzo
ph/Lgp5rdvy+M0+DEHUwnKS8Lp6XmJpb76YltB+9kRDGbvpNOb66syH+p6qTAmwt
qthTY4BDKHuRUNV2mveuFCBU9vJklAI9xByjfwajtoqXOB6jiyeQ2v3+sEpQsmMn
GYgWV7vuVz+vXGvFYlrUkscFjwOC63lNaoxvzrU5TA2H8cG9NNWmRpgMCNAvlrZA
2iigaGfc0QNbO+GLboIDb/0bj+lD+lj2Sg59QA6Ip37lyuDag0a+dZBQkF6bUVYq
IdepB+u0O6tG3F6MMKlkIGltZa+W5F2jeuK0xBfANYVP/47W8dWqpLxMVU1HTDbG
sneqoDU1XJF4waaLTpEwClvmriPR1r/tV2mkgcO4SccS+wRUAQ3g2PjJExupCHOW
JxUxumek5FFP6lJqHtd7ptqaRxpDLLpGaEZohf8tHSi7dbEdkL7iJMQ+0k6jKcEN
ozpKks1Bs8Ea64gikp/b3hT4MjnieHmR7N6NpsQylYI/OuppCi5zTWSH66+CWQ/c
8ulfspkaYqbDIs7YBZDl5zWJ64MmT86Cw+ySZ8ZE2iNIe1IZW+my5DbQdWvqSFie
7WYt8MXBXoKCcRMlFJiWxShiHeH/0hk3Id1iSdbNwU8MMO27opoFuAPD3P1QqISG
8PMVe+kfy12/binPm0D3B5teoY9ofWOD8xD2cZ6KS96OlL8AXKhFmVBl4/2rFoTu
8P7VkWwUItMBvcyicxuWkOFmOR4kVhYlKP2WIaByxge77Z7WCyRvJXIfJJXA8Jzv
DI/KNlny+tgzTZFi7HuYJxpJQPbbuz8Don7+dKIXIDnQh9QzWABnVEKxTiH1ZMGV
9c2PM9QQDAWdrCInNDYS2oqpTnaKF2q/4YS4MVocj3Mv8rgmArDDADKHoLgHdLqn
Vr+8eL4D9F5eZcS289BGhWSAVLwjL0zgy1VakISygUoMPgwOz0PbqIIjS9zRBZSm
jRYDAPZTOHVYZ509c/8JklEK4AIwUSmjXfuuxRJ+HmR4mYjcDiesHsr4Q/9Zv+7c
GDyzqSKYE+HYmvlrZAk37Uz+tke/Vx/XeZMbl9e8w+OYlMRYdIdJSZNw+QCJAFnq
LSS6aJDG9KlaV1jLPo/gmTyjnn7liuWvTDDzU1/NwmPbYGsAz9LTI3sYq2fEAExf
sbTXagUEePwU9LNra0wp1D55sJsi7GGqaLXUHjPglLOh17NHOqtsY1Dk5ueLE5Lh
nOPrbQ9iIAYHO4SHdmT925IlLyaUXc7Wa4LMZRN6WG5P+J2leacQnwzMCHNSJiY0
tob12o5u/C182ysEjmdLpyE7QEWAV80HOunimIPSbnpfDyBenQsISngBsH5yciTp
n3/hvNuizsPRR3NnVaWII1I85m3Vrs+VMFN6X/hjZ0sCvG5J0xjeJ0Q3RrnBIeLX
0dPmDWpwhM1SsRGd6ZxG0xS11W834G2XX8nLsT2QmXU3R9cir1prx/KtpiBVBA3w
07UlOQ0iBAnlVTuPTVI83b84iNPMUHmkO30IOLn/rL4Z+3tNQPT5/xCBcXlPYPYn
Zx4WAGAbLCPQ/U3CYhatuQMlCYb1URcyVkGBBr7uTOMhcTXfVcXb85kdW5qMr0sU
TFD0lwuc6tSBJEJTB8mdwU5658H1b69vZxl2HOFkm/+OdE1NkgZVITpEBYzqbhr3
eh9ekmUpCdEGU6nEyFYd2yqq0HR9FnMchz+5Wuzp2u4xAKFpVpyVrFJ2G3eAMHuV
fX9FWkXgXWzd+ct8cnLg7G3CeJGFqIhwtoLYMwSxuO01KYrcjzKvboifxE4usHDe
xLT+7EyCJN8GddJo7bqmVcXUvPJpRRv8Mc0G8u30U3309QvPBrlYYAWbPELUuJ0T
kdiOXy8/FN4Zn/Qki+1hhRdNIG4QQmOBlUFNzdrINxPILffaC45aUdLtJjDmFPsX
b6e4wOfj+g3GPmPXIe+q4c9FOL/Z3Ghm+3uQx1ebHBIWaZ1dWFjuNoRBZk1e5EL7
OX8bkMA0l2VRSVMi7CmcInaphSiJ6xTCk2n+ibodBQwr6xqqZdyc3eWWjGhh221i
HDQt7mdPfY/nY5QoOaFdR8xgRJLTGFkZc/BqA/6DP0WAUtKmD0UNmPjKWNav232P
uRBbi0OMyJRNRmyxLInLTlZH5r72U0GGQzm5m8jYoXPsqZHKllEtp1VjjLPXv8p4
FG06E+frZ1iEWzXu4d+lL0PzMJNLYkwLoy/Yw15YzmoLvLLWU7HikG+7yZ7hDB9a
oGvnOXfWhey/WyUTPdzZ2tSsWjj3MUMcKPryru3tFE5dxCkWqamONmqB/ddF36On
9vdJB96CQW2dZZ93zUGffylXC48O6Hx87Dl4yv4LA8c+fCI8De5oWoZm/KuVAgI5
YE9YM7fd/dyVvAsb4SnXsUjmHa9O6t+IQoOGllrRU/QFM3PRgYi1hmaO4bnZFEl1
8OWNT7pVE6DFZTUblmxJyXui2B+WLUHh6J6J6eazOfG4qOXwlONU/oIn7dkarsdq
SvTNbLUKyLsifXuDO5LRSDOezCuvamSrCsOWBb/JMSNJfWQpOxGZdFU7bo4E3fgX
WNmIhXdfuUnxAlqmmHyrognKt+J5rcn/mvJRDG6/FD6oRTMnUGY/mMQnMvRWrxkV
ickxsMwSITEPJ11RpPpHmV6Tuh75Qa6NRm+Bwpaj4sce98R5yDTGiPWVf1hQPphW
dnpC+sgNeYYZXcDwGw74qIGB7tds2k316E46XfBXRZmBRS4B7YElw6trDw5MyfVL
94RH90hopDhT+IJtOpTi1FFFCll/amNPEKlwDUsgwrEJMGxWVESDhIzeQJNsEM1E
FFkDEk/sKVm8raZB2I7PBQDgkrEWcYf9edgg3gKDosYNtkP+IEttJ7Qgu0ZCAKkU
mhnqsVB414GvOkgc0kM3TrKqnieABPmvjQayrevaYSu7vbWfszhtTU2Mly/XFqbi
DPU8fftu2HGvKKEICtyyojqNTb+BXenvf3+hgV3CqKcIZCZaBJ4kSIA/utrFOssd
K2lBtU+ZBSIepz0YJdPeO5r1CtEg7AjPoMgMHAbF5XLL2pEz/8jVcskHIfPpgOPs
F4wKcYzK6/fT4Vh1SS8AsEax2M/yynNOxAJMIfe4YmprHtaRnQL7fKxmh4M3oMa7
I81fbdHqwad/dbRG3dgrhzDD7jyikmLgH899atN7pVdf9YsVMsCGVUocWjfD+lHp
oZpJC0pSGKRs7YEW+Rtlyk7xubYNy7OXqmj/cJ4EI5PGF6+nHQzLkAFq8cbNex6p
+TDNWKSDeZvDVxIY6/KWr4DZ++luvUzoMkEZvykcBP6pmPX2KFrD+5G3pZXGHfLD
w/pcaUW2qPPbsB9EgCE7X2VnV5s1Iml8k9Wfy+ahW7HktrfFMUSLQ0NCoQgPXBTv
xhFjVMmLGN56390PtFUNeFf6HutPQjKNlRiuz2aVBdH0qaYGFQOpawQH26awvwGH
f7t8rSzPrONkcZxv2M2k4zrTOb19ABIn41Mnf4JZUtL+hWAtalRtLTWUdEWVo02E
HaDAJTFBG5CERBfEn5mQoT0GnSX5ANa17osUt7Zd1Lk7/qsfhw32jm73rHWTevZT
q3IgIKiMOkgMLUpzz6KXDnIVgEUIxRxtm1HndivsA5H2YOHebImEjywS6VTeUcaR
f8zVrag43pt0nSuP8DiF1e8pX1woNnGNRh0DVo5J0lJTpXwU4rH+YpyQ/BSO/QVR
RvV9zWgLhm/8NHhjL3nmViadPlnIcc7rwv771m0Kcn5D4uO6J/NN/de4wD3ZsA/n
g+iQJa6X60hjenczqAByvg3SYSqmKSgDTcWdDpBpRjDv+SNeb+13wsWc6ZC055tZ
YIp2e4bSFc4+IkK5qxj2dQrCIKD0E593Lj8TwlTBirY6YExppz8a2FqLfrXYDNsC
+lcK9uVNgRxrxxE2CgRGgAilZ244VjFhRvgsJIEsVq2dEZ30iO59m6laWHYju5tT
FjtFwkmfd6ndQgObqk69CFRQdplFVOXow3O30z5W795cdBCeeKQzKApzZo9SqaCx
Jq9v1M50Kv1n5ewYxJ1RmwxT4zh8l9oCxfdkiR3t/pxsz6sQp+x0qrihODb08QJB
N3TiyLSzO3LDhYr/ySr7nZ2dI6mAcgOBFcJl9vgZ6HYUpyoG0jZ4AJs1XEzvvcFm
5sJsRNLJwK/YEy5yvFyfA6FpOU2Z/lA2IQXU0s810GzARmR3BaECmTy1xWS4cuwV
0wMuZ11MDSE+TKsSOnyl6p8B6kUZSWgsaxIF40p+f2kplcytAAUREkG8jl0BBQ6z
RYvSiVQYOCwEYOzHGuBKN4QHkpppz5NqQOGXae5rk9sRbo3ArDSRVFkRd3zSSUTp
3MOMWC0WwcWqYs3EXU8PVGw8A8mkbkUZ9wCAqEqEO+/iSJ/k22NJDdVXqOFNcmEN
+KpTm1/KAuopOLzDWPt9cbUoC2/iSTfM7jYMWo6kIRuaZ5H8M2KvTP7GBMe70Uj5
K3QxMsFtgV2vUdNn2KjK6ajK+wvrEBJv8p5hcTh2qnDQmWdWYcZhRE/DinvE4ICK
Mf+iK6g9rT1Yn6I6Zt3E0F+6vH1Eiw49mwsO8UcxRYLTOppLgAumXF35ul4l5eiX
Mrt53tGK0iK1ZOB8l2BPF0EcixvVaPAAnDIXeX++X+jlP7nzKW283zgh53Ikrfxa
O93oazh+Ocm9FGfpcsmGMKG+HvlGyrc04USsgDwB7hQsvhunWzergqACI37kWt6H
cBUrpASFaC1FIjtW8DeWJCFeW+ByXbiZevTw5ThvUafDd0c0g5QWaLLuuEHnS/Hr
HYAd5Yv9SGAksmAkX7hi1d3iY2u4GbHhd2Vf3xWqEmEDjLh24RYp4tKkd8FTaLfo
DIhafQZREV/B0xBJF6aFqETQ/tYRhZbr+lmyPm1QSO3MN+DbqsI27p0Y2nRkrlWn
BJX2STdrCzHfx2vZBWwEeZH4CE9IihBeV0Mi2qJfZvr+NbT+zNT+HtuElr/EcvQT
k7LuSlUBVDPtB2aOE0Cu0YWAWJJWkO46ecl/n50SvrEQu8gmx5QrFpLW87V3Ck1y
Efl22B1iLPtgb3tf2uPe8G2KTpvGapBdlhnsCR5nfcslreg4XYaZLbLgQGmvd2PB
2vCY06540fKFvVtN/duEemiwydwkSqJcRnJ+REvkrKvXOt16Xrgxn53g1OyosUt5
5cb3u4zSmpGV+4NS6lx/KIPfqpLyWU6j2dD3FbHXI50cTZdH3Njl/67XN59mii0U
YxgY0J4KVMw1Q3+9lbL61wEgZ4oXUSNTIQfYB72KsjC7WKfiAKG1yKAxm46h8icR
exRfekAuW/k676H0Djsnx9FEGZ4P40ZUJTIjuPfTLD/e97CvrzrVj6puma0+elTO
4ChO7KR8Sy8g4OzhwEEJOf2uDmfTpR/USbJv6KNzNN7VflSP98Wn5jTTYWJzEaTg
/u+U3Uxo+/GioDzwrYCLjC67PBKGRZeI+MyF8EzUSGezpNasHekJywN0XcNoHKao
eN0CXL5iF5Z2BJfFtUK3B9jQhIbWnF/HBzinUnp4qwJesxHiRt09H5xsdNXgRExx
d7BBubgu7Ktq8uM/IoVy4H7GXNWgaA+0DhWoR5/CvS0qKfQovQNCpjJ0JLSh9YEB
bfiCUsYgZjPWiiV+pCd5BMfUHVGbXMPvn3FLYBFq04zFCNrjCyxE4vbW1eveN58w
c/HeJq1yeSaFOAmdWSvgiqYWFIdST06fZIt7ucPsQ76lBI++zTpZ6DbFX53IHNBU
4Wt/6+6r43iC8MIpY1ySJMAeso0QxTF4/xPue1JtcCFYC2g47H0piQAVKXLP5jcw
6DeRWE5bNbWwuLubUN8LdwvFQsEcijT23VF3SgLSqhI0F0HULyLCpTBguk2Rns5p
o0ZErg7Lc8W2s5Pxl9h/dtbUpJ+PmZh6a4+ADL4wg8juVwPIb1ab5arDOcDeKeD8
PNuuoA0qF9aJc8JNtotRhfHYZyfvBf/DhZ8BYBuKz15Ir9mVu40agCiFaXNn5odB
wmn2CgahNhuxwCm81adKZ7CLSoilWMZgoNP+4gOln4gw8z7nMGCMnx0kGvrVro0L
pwhflycAL15AkOTnLJ6K0KU/Z2BF+lwD7pcaKBneX/FSoNS/lNODbjxwbKjL5kHO
3feXNM5Ez28U7IPnKP1drWpiKPYEEuM7WGf/vs/YnLpq0TLD71TviM7sbjlDKVwL
hdyoGDz+jyEAbI3JQzktDAlgWZJvuVe1gk2Wh95/caXAgA5yp+4FUXz4bCGG+Li+
sH0fj7w6idNaaNdZK3NC0GwJNnbO0QPhigyxUdkI43mmlTZYpaTC/C9J8EjNCTfu
QoEBC0Pa9RRhU7zmj5rixTL8uSLn57mDy0CkWPjACYw3gUPpTiJhLyxf6ZFFsbW/
PBvAUjFWi9k1FUxpJDWLTXDiGF3Qa3GYvGKMP46/+ttk9eZ/09dQ0WDTdiqC+4nb
1FMQJcf+O6woa4NxlkubSkRd3lwODF1mHd4sorFYrAx2/vXWhpaQwj6La6y7ZtO2
dMr+b6M2X+E5ju29MpLWT1bHRVtbCYhGO75Y4PwfToWy8VrDmykSLrzSw5y2Y+Sf
W0ZSxqAN384gE3r0RcimBcqW7T9K028VKmqR3IVRkH+p7HlePvjAE2raSJUEHmn2
0Dbg2gd0noHUd2cfTKhx5gzortY6/kNU5iWgQmCwR6gCPD5h84nKAWPZT7TxD8Cl
aNQYty0cQjLrCGqBDxOW0ZAPDutoIJJEmxLko7iukvciAnD+q259fl1uL7/qT1Zv
bI/5xTZIHoGbiT7P5TJBDlbp1WIHV5feOytIIw9MtKMESVFDwMa4GH8Q+crNjAlZ
FOwzcTtWgrqjctcCy9nWNe6wlyyIaQ3BNKEnJqFxqvIhlGkrIIPBP7gCanOql894
TOH84bqZocvZKL7IMsbC8EMXwNCaPEWw1gxK/+fa6vDvUs8uRQOG6nPjn9/MtHoU
WhoyrTkoxl9cd5X66Ho4Kp4B7TOj6hAXOFCgPE6+lb4YsOlHWSMVyJE7de2DKNAf
HtQIJ4b0re9rG6a907MNIkjD1Wr2ub1EkpmSS9BtzOUU9uzuwgQwJBfRCvCm4LrY
BeDlt6Hi22pomFKjSKqE9brk7I+1LoEyyGttsKldSTCUUgTlBU2UG/0DHDBeFkW8
5ApaY3KgHRfrobth2fVfwaeyJYGrKzvQ+v4/WRcRHqD8ZE4vvXdYSILXumyrFJW0
LDSSv9H7Va+u9qO8BAyT1mttYtTusH40EXW3qR+1R1qyTck9OouJE+Qt07+dDzPZ
EzdVUv8vDtn0G7s7o7kjj8D0Ug2hk/nM1CgfaJvr+L9Jgs3/+2h4/mYZgve/jdDE
P99TuyYDHgKRD/0wHN5VmwM86S04anzE6nZ/dFf13HeoqenkbFVoPufBMuiWVQOe
nbk3LzVLa0gm9cwvJczLWOTqKzRtzVHPymGKZDCr4B9VUIIrFME06bjKJscL7CH4
YDsGs+L6aVZQ2EVJictYKjWcqP6Gq9xW0symL2032BG2dg4l/ZllCUnHDZI30M8U
aUBC6PT2bdrZnu3SEvZJlOQeXFfmeLJO0gk8nEys7h3bELl9HH9mnusprOhj/rWJ
QJbh6HsRPcqwl/5MGxDDNeSJaIGFn2U6MgcEEM4Eo2WEe0Ol/z5VrxPd5oBIGC9n
nxlez3bqCI3vjuSsDi2OqWK+Z9nrjCADqO0jU21ead5i+8dfnLrtllvDe8zmBQ72
AmUChy6qvqSOZ2AXieTPw+TAyXxMg6rStQTVPDKAOyV0gL3WLOk4mpfpwtSPKhNd
dBWW5hqKlpk7rGkwwU/VXZVNnNOB//JqAROHrU34xRLjy9MIW7Bg5uI889HHULIA
ck5WRpJ/qnY4H9jHbO+y4Cta22UF6LVhyquiMdMD16u7Yyyrpjrb8feD5OgUPj3K
v4h/JvrL+SRqObhTPbhk1DpMVr1ddlRGtKWcA0KKn6DnoDSYzZn5Z9j9xIBxDXQ+
rldbreDXBzB65I5s4mp/emDGscw0jKiUKj39d++OhJb3r04jD7CUSQS64MHFxD8u
g75Azxm08rLvC7xb40+DN/IPmm6i+FPkU97LmnX3pHmppWyeSDUMyEz/vCGhW0jl
feV6gBBM9u0SypQrkB55PRk9aAhnvak8wTWlxeukf6u9WJQfbqcM4rC++qzl9IEQ
Jexd1eMNYyj4QNzdU2kzEELZhr07AtZnkUzd10/B3wSBlQdmD7ThHYgHC7WKPSLk
kKZAagTwhzNtQ++gm3sifRg6qG/9HrZaXerFBcB7nA5aE5aJ9o3+/VUHaxO0DeEv
N4Q8H6SFfqEuqfCK8CLrtbria9ayjMifePlFk+E1+YjHP7uWGHY6RcwPTgjsijV/
pM6KLcl642QpeA+pxkB6tEGI0EjPJMJYv4ixE9a7c/T+nfZdYdRy/tMVvElE0w/F
mL/u4B9e7RrGQFZUqLObRO1XZWf0b+V6XRQkVP9yVAr/Z4lwwNtEPXUHWmbzk/GQ
B14EzkVMaJVI+yWAHVAzMwLHyxN/Gz/3Psf6IT5hMcs5FwZ27kWScJv2ddMvdOBn
MXXWnpSZZXqHp6CaxNITqbCLQNZRKfdNIHHq4U0BxK1EFyJ7ayrH1tM6ogXTKvgO
s/0JjbAACsxanodIbgevQ3FoMMJfnBMKGnjCbv7zcJxBOrUGbUuwzK1vBJu6r2Kj
tb7HChR2i3E+SJ/YvcE3GFPxgArL5I+elmv2S+m3n6VrkOi1j0UgZU+dwuUdIPP1
Z78RNf/8qMFzFwe+z0BobD1zuWjy2zg8Y5HC9s6WsoKxs5F84EQJ0cwvddax4Hqx
Mx7RuifNE9MnFUAHTStXH/Ja2PNF8CJtgo6jRs8Uk/0k9pVCCuixaL+K7PcvhSgD
aoEgE4scHBaTSY7GyWDFJDI9hMXCqSHf2rodyzY8BwxAJEz0R7u+OagemTVVG/nq
WCe8xu2lQiUkcmRTJExj8xdQoNTEu3CsmXjMbKyzaLzn8Ym70Wdc5V35C56VZ94n
pKeZfmrCkaPab/D+wxoXtSsmKUDE/glnkV8BabsvJRiCWgBbMvbVx3ctp/1aKWvF
sUAIo4P+9K/HkpUuskdpvXDdwY9sj6kQ7tvZa2AqqZRUSs/zC9I/31z0L8f5iWoT
gOuxpd1svqJlIhU4OLIHyvVob/5EF61v/wsOP5UESZH1A+yWgb4+0gV03ZA0NN0i
LXIqNQ0Fb5WrxpeFmVfvsHAuWuRDreOI7xlTKjD9hUNtaPcTHsBlWcwwXdvosvAs
/D0GDW54Ekv3JGnn/siUvcgsHFUTm6Dz+kEjDuVteL632CCspOYdoyrJfF/Mlh6q
bVKfJCCOWF8ItTMlFMYvrliN0bHLq/kdrPOIyXi54ov0G3YD0RXXAmgde3aHBz8m
GfbzyiBL2oWTBYasVbfh314SH8gT+uEQxUDn8BxwHSVSdOcvgyLZfIl5/hfm9sKq
YrHJO+ueZT/f0JhqYd583W69cusUcRX1oEthu7Si4tUNazn0muuVsfxhrtMrkdHr
3H5gcL2TzslwC4r21HE005H6QvKSSzNCgcFixCpoW0z8mFaP9XypOlzYIfbGdGcw
EG+zM8R+Ic3Oebm9DPA2XH2BzqT6IQgeCw2NCDgzrnO/PiWgS5j41JwLWKgmiA33
tAboYrQVvy3l/9wKhhuoiu2h/FrmS8BHGwEt/OR8S+R69es5Y3fRescvQhPyQAiW
UqKSJJWD4/M3e9UwO+cdY6qEVk5hsOk/rGTSpSvXoS2dATLohfN7NV7i5+0oVhEq
/T4S8COwow/bE578TnVwyos2fsIAZyg5k23hI42urjzBCjzjwBesEyI7hCCyWFoM
bqpw+7rBr9AqD0Ik5vaSfILrDFBLQdNcpDRuOvkPKPEoBuJjB8j8PBH4UU+gmo8v
ZXqK+EsXP66OjHUUoCO9Xx4v4WhX2Xwiap4M6sFbd6jrf5vT0FDDe8EXW3g3FfaK
hd9BiQFoOQqN2WZwiVCjVr5+2YODXePWHjvHDU+wXVj7Anja4f/9VGjobMikv4Lq
ITLjhyrCqHLXUpdeFAJqQhzC983yrxTCe5oNcim0IXLn1DHP652qBx50HbvrCYjz
pt//I5BXKkUJJ0Bw0j86pn58MoRcMFcmYoLzfgwfZML6TtB05PUWTOAAuCvB4KKX
RXU2+4nWBBPDOrB2qyqj/HVh5tt7EmNieDXaPm8vovE7vti25rX9mCpYXnw+JiWW
Ox8/0yh+XcFDzOogxhDiCwU9KbZcNiaFhB+ad/Rfnd2fG4v1rANT31sy79qyZ6bD
KHWeCzgqT2Qok549Smqu5mAkiYM2seTvmNItz04EZse4mWuv0UuD1pONHk2CKger
xS97kfza3Iu1u58DasvSYdrwA8fFSpTNM0vvnnKRW1Da0qUJS9uX9HOOlCuwCuEW
rtYaOrznKt8w93GS6mKKlBYW0Pf6dBku/W83ytdHGmR+10DxM9bXfAMD7v/bisbu
8uXSt2oxGU5VCpvlJ/cudxAC/5P62gOldIsqw2nvB9CufTTOdNuTi1D1rm+Q4ZES
9V7us4knM58KkJByfNCTMwZiE/bDdX/BtqjO+7vlViYIFrkAmQ9NHWrXIJxJkHkp
lsG3UfyBjQmYqStZSfAaxcy9Qw835Be/HhsIXVw/74tMMj6jazs324Vzbi1In7md
HBj3LqBnyc/Xhaknj4k60FRIUaKaRsuTrDQ28OE1tlESbpZkYdYm6uiqpbqNbHvr
SjUl5N524JVvBXHdL2UIYdRWLW4hGzNaxW2n4oGx0slxKsLd+hgauhaVLuzSeXfD
4aJ1S1VJdnfQi+yCdYhWYiFsUe7hGF1LXw5LrBxiHnmnYAJ3I91hWgmZh7IwA/2K
jEsF2KSPhX4U+fEnSSjLclxRKxxWt29DubxSmB6KBRFqj99LUCRJjUZLjLpAwMCT
rYxGg4JeIl4yHnLofBsh45Hf9ILFIkm6rPnv3XJoMoKKXj28kihMG8rH26wZYaBS
KrOegHpYYhH/wniFlpmLpPoC+rzIhnxoECHRtr9QpDlO1P8RneBTKHHgLQ5FsIfp
RlQTMubMBQ6eTKgZ5wldQ4hnREdv1nuj3YZIZsGkBLOaUwvJrclVMGpHuSqO/eRQ
QY/HcU0XID3FpDPlFz4qvF+sS4JJGoL0uKKw1q/LQKi0h+kCFAxpGgzD/5iJqVbE
TBV50bnv0XTuWIZZ/CXck11K0z1ryHjeL888KD+Gn5/Wtd5VF+aHVe+bmltCJyr4
NVThtOLyikII6vD6JI2al32Z2NcDOENuubTvo8X9dW9zLKHT3Jdof5Mx3UcAk8sR
/8hQ5LczarMxUnUM8i+/R2LSywi7xAvZs0f/fkFlTbSoQs/pAcZV4XfSPXJ+ZB+t
5nUOAvpAhj+ac71feOerlrNTQGyBNVUa4RpGdeBp4SduogTz4kzXMKqpP1DXnJwE
jtc0EhIqdDeoW17ZBFo/YZae3q0J30o4mU0VCL0DGG9zllgIN5aZ70hV04YBbsmd
GJUZEg9sAOYnISY5OABkd7nDs2tu59SQc9ZyzboRrGMQEpQNYHu9AHfm/W+qolXq
OBSPca1n1kfJGXX/ptLJaPFg5ddibkBU6IvT96XACWBicqISWidvjKgguhvr/mLz
X08aH178hw2uaWTnJqonTGuX7vdB253Lnr201iK+IRFdo0XOXf7fkKqagqhgqABG
x52nBUBNfTTSkaFhIOB/xRPkw3lykitMGylFxyJpOaCpGd5QQgOH5V3OtG2KNRrV
lvMJypRXWBjxdy+qnm5xWU584392p/QKshgIrfZVKII22PQG0XsLXQp32E3QCp0f
atZKbIDOdnCiutsu7xPGv2nFpCccGZ5aQWcc/saqjv0+QbRpbx+LJ+oW0rPGavMP
+FCDdzKS8dNWwgDGg2cbZKOiNNM7MjT8wi3KW/X2L5UYfFWBfQEmiisxi7hVaNY9
Lv3VCNDlZwlbkU4NTblsdaxMhgrKc0x3Avli9XtVzxdIQcCO8qmjF5VumJEakvsP
A/ieBTqVgQWIKyDNL0UxjCMoaHme1smoieOmI6PPz9Q3r7V+bvUqFDDHiJ+1GZ6Q
l37xGWpLSsR0FzhEAzfcXxiNnlVkO237j4loHIgMk0qsOn52erVFFlwLSazgtKYK
RdR7wkI6kcCj6/wP7l4sJTe34Ro7z0m+aOq8jVutpwYR1ERMLa2XTBcrfdgsx2op
9XVeWvjCARRMCfMmkWCotri2oj2vGD9kzfbbnkMPDcoWXR2JkRsCEQStVEc1ZOtH
GYWwC1dg3lf2eidlSeYzPbn33kk4I14JThKOPYHY65uizjlfNDTahhefhHgIFtPS
dLFNhuJvEVX4Ie9IvdZX/G8J9yNliBWqW22Nc6dmbGvPqv0HkFuezPi/jxToyuBx
vs/9sFdZweieMZcmjQ5O96A8nm1jJkbr4wvoRk9mv+ln3Ii1R4XtIrGbvboKVzgN
vz3RGN0YGX5cRYxPIGRmqI9+wHeucS7xpyW/IBxa5PnQceukaypTJ8QlFHE24b88
5oTcqUfIxuJgXXNyWNT6NviR/MMItPOtqRoRG2FzQpO4M5tsioCWppQtIp0U6Wpw
cL/kCL+61ENFLJIBuQnQ5YWIwkGK6wC46tpEC6MXtKZUzHKPW45Jb4uw2V+6G3pq
Ge1upt1883IWuWrLoJTtTHnuL1jbWYtET6AOs00iJuTa/R8WZtOK2FLhXsi3PqtY
aT63JLgQZR3x2F2fj51fIoGdkuhbMjGjMxsOq/l3/E+VudWvy5TmUdYFGGvr2huw
ZBkWH2frTv2KLOLYogMUXbfokYX9oni2VdsCsDEPtNJysYsv07gr5tI21h9g3Ams
Lb+MnmR3XLsKmaOoTD9X78u84TXlwXkm+Daxl7zWhKe9X2G7X8K+PF7utc81oXAV
Dj/M7PIL5UzpDvWKvc2n4sRXCy6f6QjcEMiiqwgH1UZazU+mA2tZSiv6sN9kstIa
OvbZGVUImwX691wFczFfWnphaY9e0cae87az9ILqlGBMvTVV5qTHVvg2dpDifLiE
I4rZZdjUUED2dEn7DDj3k/5rysqvSLU+9tHH10VuCDxVRyY/rh1dC2lAH6wdh0A8
7olyF81l41D5xHdZb8hWL7Rne2TOsmhzkCNXzFmABKSFPAVVOBvSNiBNQ0Zlmu8z
dq0Y6rYh4jY3flLpEUXH03N/jjO6z4IobzXyFq7DcbYQPhwICikoYKtat4wFsjni
/zehK13btfQib1g0pbbWRxjbBSiRA+GCY6d6G47+KH+HKpJDvHq0hDGYQoRR/Zbc
T/fXU7+/3l36Wv7fyMcY0Jh2jcE67iKoMT3M0cvDnIPZCQ2iPxcaO3ZIhyW1ifzs
fQeD1NYH/+wmg3fD5kvfR7NZhe9W96suPur1qh5NPEa42ena3f5ZHmZQPEwLUnld
kmi4kf48wHvgiQoZRe3hI2X3hgBPwwrWDttCRyi5liCNJb1jilTRwrCTP3SXaqHS
EbECmaPDJpOdXWVZM+z/FNNW/g7SCdBpYQGaQBptIiinCbLZtJIjIZQ+EJg01l5k
2i4xx6dCs74629dkMVlYCafNcdGlbAmmMUDm/lNQ42JFZF6+hdILRqApk9npFggI
881bN6fqYebrxYHPWmTLYemcuY4uQphbpsToFn48tEooDS9v1FcvX3COFf7ijvrN
wa0CUikzmTpXlSriAJHCAzaAlWNbRAsz5k12EjPfEFHgsRX6TYPwoSDS8zyObpMj
V5//VRxJeoZAHGkOVqmn+G38MYpmScqhev2A31NrHRXmSfQH8rEIb4VOGqIwKQiY
ZtWwzzNVclUA8uUnZnyJU8VTMFf3VV8MuTS22AfT42jjOdeEa+RHEej8UEMV4O6Y
ikr7YZRSVR/s02enZ7mU4UJV4EfCE57yZzvwEVeEwPH+ILe0JhbuhB4UzCI64XUa
M/SFqFYE1Jp7GAlVLIYbUi8VXxRUW/MQanYHzzUkC5yanhE2fi7xkUJ+NB3ChNaq
DWhHj1JfWT4+Xl3IM4q2bay5li+jHzDjTWztWBH3a+MawdGOmXKm9CAGcDFHl+V2
ySRKJGsC1MQoBYV4FaU15BQ6lhkn6anuOUDEcApDwAncKnyxpBjuCwgstz5A7l1c
suTfEJHccHbiniz/0B2qaQbpMDqNNopd1+PV8qgXKwGAhSCwO6oFLZS5evT95DaY
HwvYRG+Ik7sHT2LzwavCEi7FLilzV4h0AWhMyxibmM9OwXbv1DSEuAaZ8JHzNBvp
5YzYm30xfrzFQtzjfOvHtk3m35kpqi8aN0Gnkn1xNIhywM1m5BCEHyigkxMymBVL
HQA4hsrThYI9RxOecBtHHCB6PBt3juEjIOz+5tbvpnWdBjwAQNEVaj8h1fAeyaDW
/kBIXeFQFvlimvA7JkiOYSdMF+4Fcj92pwdsAjCzhBtKNgjggD28y17i99So+4v0
3rJwob42pD36edzDiMI1G7vWd4PA+Y1WfwB3WyBovdj6mkZLKM2aO4Y2t4W0IaA2
knj8NLKRQMC5PkFADtn2gY6/LjCOapcTUY1/Q8VB/+/U84is34/XqgClVPxoBWp0
0O4MUmErpPmEXO8QMRLqqAV16n3OjwGTZvQqTMaQdFHZ+oobGhxgzVCl5SeVnvzJ
D/kTWIBBEQaG8lmvZYCRACaMdIV76OuVep+pPz8rwvEzdaqzKt5v9tyXsPN27o7e
WO1B2CGyS2F50DSaTm9LsGaUrjosdXfAnpgdCw7rwgLZ6yOo/ilEUGLpNdgZiYUA
KsSeGnTZq9+TeSWh1y6kCvjp7C6x9Nrahh411VM5cTbt63rteuSt5KFb06IM61At
X3OSBfr1GfYbh8VWIx8jwXaCWUxb+aG28XlDp07yJ9Rh6DFjGIDEkMvkI3JJdhAg
qCCfvJ1cWKwJk6K6W41QOjjJhqlfCfyMwAJxSkcPfBS6+dQMGEREvG3f2msz5LMW
kSBSNaeEEhvzl5XYhj6HpRoQZnAPbZnnyynzUJZt6dlDBUOV4qtTDqNi0mA9eWRE
FUoYPUiUkBZN1nrk/mNqCBSmnSEImzGm1xEnPF1UpFbMxennq4GMbVEqSXemzGtk
RRipvxrsk4ejLXlzJkdkmzqzb+l3D5AAcw63qpYKFbsOaF66sk2Z96GISedAIaDd
d5gCpjn2GBTf7evgJCXsEl05KV1C4Fgptw02pe/qgKwJlxHN+6JIjptpD03yyefv
NDdynXzfjPkHDmHJRDXENfUucsSWDChjzyCO5hsUSB/cD4uWARKhEnp05fjj00wn
k0cc6V1xU/3L/0M5ksQSGTX94WSbO3uNXE571LWEOnLcGEdGDGnUZczBEa4vfgEn
/FTxXNUXD6HbOS9vs3YXRdNbbqTVxlE9ZCT7m1fxAz4OXwbjRH+dNJ5rp8O8ohbA
X1OToT9zpfCz+/snWWK7ylHgSZGKBspbz2LYt3bIvWzgwin4szQfa+ElWXDax2zS
LwdMDvJAf7X6lF0vie6O8Hus/XumL7dXiyXnXt95RGoNWXz2CR1kBQrOlqAvJdBc
GoPF/TtgQjS48VZjacNaWtv0PEtt8On6wglyJYxsQLFHesoMT/BCU7GNmdFZFa2C
w149PQ6KWMWx//wSoq3/AoxIjZszAoRigDM5was71Naxj+Daf5D5Od88MJoXN2pg
Pf1CR3beEHWor9bUkSY0lxRoQ5wkvxCoWxhRjk1+CEdSyFQazXhiVrVnKRwIXdv2
9CB0nruEGo9fobvtM5tz0LfKBxVzeTLd6oF9rdzh6MPzQPAaWouqfooV3lngZlU5
DFUS/8JBXuHNTnEpkx7Qo+fRk+QibaYqaOe4KJRzQ7WfBFXXlmY5cQusAJx9Pg9y
heq5Ch0MWhGy3LkgGkECfLu9W5rRyvGKFiTz3pkI1L3c5+T3nrLlFbxC4NF4C0V1
eZu9EVsh18/bO6zHQnt4Z2EoRofMoGauSBWROP+jfsn5uSO7OmvipHW2wjvBNeKj
3JW3KLDu8tf1s3WZ2Evc3jZIbiG9KSTndCJucUewFjAnXr0DSws6ofRPwRvzwbcU
Ye2EWbdT5pPLQ7mNevE1/8De9pgQFPWijjCcRJokH5BAjgKT74bUyN++sYolVQL/
N5JDGXDQbIKaL5nFc6kiDviC/JxC5+98lA3mKWDh9N3O2dv6Wb1mhjG8eP+TUECp
uzREFNsZJYa89RG3eqFQOVVAs+wMMBFfZYP748Ql27Hx1Xmh/IsWYU43vfzpIRY7
lEGHTYdFrs32FnvTRPO7tHa32yYAkf/U7h/1HB612OFtTqI5il93UDr7tYy3kXd+
+I9JuvaMCWjhQJ2r4lQFC3sHiRyoU+rtU+/13DVeDFy4frzJ29gJ7bm5mkERbOer
BCT/KAeznE9bE4e+HaQ+VNJ7M8yISw+g0fYUUGqoCrrr97mbTWL22TqPwGfsMNa5
VXP9QJQ2gfnxlbNc+96fK21NhRKXYmJ1ngZsNdWeW88/oFmt/IBxXT88tJnY9ESz
ld/gnuYssrVWvYhjXiy6M0ROz/2VG/Kl9i7kwW5/XMCmRxzxF2IHe9eZTCpX43wV
74vZE3tLaxw06AjlP8KDHRI2C0gih8iZZOev4HtJl8GFAib+q+gY83AGTvhvAr4V
2TqgUVmWTHGIf4K/6tVH/86YycqcXsJdEhqO7C1Vwilh+YnX34g+Hor6c0Vi+vsf
X9zxI/0I3HTY1YGVDUndYqMKU6sGW5nfuwtGYxeVFMPPsiLmeZad9/4Qh4/0mA5+
PYOFK+iJAiNKZErkTQbTN83c1c0a697k4ps90SrI/CUPnqj/COot9Ut7kYM1C7/W
k5iONbeJNPpt0r8Y/LPmOr9U/+BotzsHT+B1/BcI9LCAkSclQVO2gfF83n2nWQlm
e/8dzJehjzVNJyVENo1mfrjhBSJUF8ajc1f9hiSBuTmKn4k5xbI7DR5pdqXKpaaP
l60T07zrellgwGvCnkf2WfStnbbeAD7Yu7ROvpkYvfNx9lc4+KA7rwwXBQyWuzOO
gWVsYCGPL3PhwA5n7SzDNxEFL2xJCwmGKZ5yoBRGJCGi9gJLRMRPar8gIIkUMpFb
HF84zep071OaKWUtnTrxZklp7NFbLh90Errjr/g+NDE8TNdWPUn1dNtKsFXTpg4g
o8IOaeDrVuvFGLvGHMOeU2sL6e2L86laHUE4DImdZ+0iHeLGx4KMXdHZ4LoDFelX
NXI40gjZjpMlsopFSbk6ATI5DuhPfjrsQuvMv2BAX/bmjJL25CEweGbLNLmrRI/Q
T3/ZjCZclSx7VlBSukLsW5BwK6QqiSLljAXgQEJXPWciAEC81mYxjbIl/rxiNOzc
+3X/RNl3BQ6a3PVkF0CfXUQgKl86Z0WaeahzAO2dW7rV3ylNGewgD38uTgiscyFf
R9C8OZn9EoTtrbjpe6iTniRYuImnMSZgjfe/+Eq2R8kw9OrdDeH8IDq+PWrMiKAa
eTD8tQIXTuLO5kX87Qi8Z/zfHKbY5kmAZObGJ+Oi/Np0tfHKi9UV8iTr3MyoIwlu
N00G5JoOZUfB7jcRNcl1f4QqYYcIu3GOulaShhNRjHQRRvd43VH9MGgcGDPdBNNW
KTnhX/eCZAWxQgWAfE7EFAYPansK5bbZcfsT24jNPp7PpZ4JKKPBFpFrLkFfR9gs
zxEhsOZoLAsTmRacvJfmcZXMvE4JCUByzZ0URCUcU6LG4TpbmBW0h2QCYrWIdcj1
0Hu3IEG/Gi5WyTLimEOUhR1Vw8zd8qd8VK1ELcHhQTMxqTcY/LkmJwy0gjOucMyA
8OG+qXDka8RebKH+FMIvmrLbrVgK5VdwxjpOH1HkKhWhDbZByGNgadiPQHcrtOjY
r3uyme+j5xSLSU2JBBfih10t0wzruVcQRqu/qCZZTHCIgpUs5/jOezs/BgJrlH6U
UqJVn0vfk815iskUj+Jvmc9o+tSIrb5AUJlciH+t7Cl51P+9kGrGOMFVwnsObiQ8
lrZc//U8n/t8Bf6siVyB0dKE38Dejp75xaVw6hAE5hRogbCTOMTg37oBPu11WXbl
SIuzhlleXrFoziihdDOLXkIcht6OIJ/0A2iErikLJIV0+yQevEnStwL64UHhq/Fl
tOGByhAUdvUdPxAN10aadkQ/Jm5YAUheD6u8AHlPEbL9gOOpT8qtykCdBSQrNReS
ThmuZ/hz3ZmVTQg32TQFIIdKQRZ+2fJXvZwZS80a/q23kQgG7FcRow8FzlIwCZF8
0B37lhd3YCCMjkxzHldeLJwLhsdT+6uucgUT+FUHL02LdasbuihaB3TBLvKaVslr
WZVJeAwf6U35oFqmTZio7DFiMjU0ySvqbL+7sAQk4ipNYpbcTJiWxX405LOfbzyq
59V7mUiC6R2gJUyLxYg5Xu0jm08+tOrJCm4MQpMQ7MCMSSDszSJo9Xi8thYA4+oM
xi83FVAvcips8eVWCNPhFGEkNLInBrQuBPYw934RBq+E91SzfeahhSDWkYCIMCxT
Fy5GJ2W6urdHtUCBBHyFFwnDrWO45vrRL1jGEzNCAMcUbG/rxZkkbxIsoIb6wCoK
Ju6ybwNkN6vCAiegDYB0Pq+XjWSY7xd3/ruqZbVG5qo1fLuJN597m68L0paIi2d1
JEH3AE4ARqzLnp6cSHHt/MV9/HlmvsHC9ADajEiG097+0401G+WxvvQB4XWAChZC
l8BJyT+we+0RnJnr7iqGRZ7YAQfkQEVu070TIyPTJM1feQttE2PMO2rVmiqJIbAh
PDxcUZY3rjQgcjXMOeRTsb62z85iuuqKjUJ6n//mQpXYjEetCoDWfHkKLTp0zYaN
z0oOeIl9HaJTTxfxbJNrdnTx2Iot0Kz67ctvgLRP2RSB88dbCum+DIl7D/H8ykRg
IvchcUvlRhuOa17rqoLRPSmp7BXP/s0CNtpOIKI1Cvv3J6ppswoD205G5g/31ubk
nKQLUE4K340pVlVNtDjJNRqo2ehtmAPAtxlFFJUF+Y1zya04Ps3/bOuHLGEpNRBL
kveyhKmtIOxC9St90BIMHBVK8WpxaXssQikNx7phymIzZgvR5WEatVP6sykDHv4u
Vdru+nLXc07tRvgtYLH16Qktt29FvKwpjSzHT8ZAZ2PoGxXPzFBfT1P2s77S+Bce
3aNkbgHanHiEv3niLutCj3z596MXQ6nWmaj6YKbZF/wF1PKq7TdASnOkorPgPZWE
bWC2k+sXS7LVJ/fiNEa/8sDkYckNGHfGXCuoIMaHzPg8pLlcI1EDZj/qv8g+2yPO
9XBdQ2f/O8hd4U4y9c2fWx4kHxSm+ZOa10HE3wpUBo7NfyUWqlAMpoa7vEAO80Fz
Tbznmo3MbyenpECQvrDRDaLY9lL32+xKi98F7WmCBXCLpFekefNOZlYJkbxeIkKb
aQYlaEakqSeLrv4TwTv9r4zaZbJ4OrqAc6VSQQMZ/zghAqHCpNEC3IcOdEAthW/r
eOdurVxDPk3MVYl9fLlDKERTXeSJSV4YrC8pe6n7M9OcK+knDp3BHIyav2TRiJq2
iVCu4Nafkeh6TMBWDHFhldLarQzSMRg/PR5pk4IFr+xDeFnBpTdsSiFMm03LnGfu
gWrKybJLw32YRlWWclgkasqcZwb+SZvCcVLBhEtnaGn4PrDMjqTGPAvBm42DezUb
WAz4uCTftQ88CGSLX+ddFHeJ8iH/W18T84vd+CfQR8EjlO2jbqd5x+hc5rNQp0GG
3ohMR3iskTuWuyLm++YevH2Iug7lPIi20XQMG6J5EWqZZDCwdimEaUuki6idTygx
fswST7wOVk+ybUyJKPRnfRFFk5GdokdZmfRcWA6D+9XmnCXadJAqv/Lm94ekWo71
FiFSmuCzm2p0Dep9FmMoUCgHoWvEHqY1ty9vtg8DpneJURka/D5yI8Lv0YI/U9Vn
RwHFzMTt1FLifSUAaXerwccuKYfXp6s8BpWFEH376w9+62fofA8Pi5t0GTi4nGsn
3otj2IzBGlPYQZzuuw5BFWe9BANWQuc9oqFowmAwDQHbF/h9ABCk1QgMoTq/2OVm
g3EaWvxbJ9kx3ED15p0TSe3sugr2DZ+ywWmvNh0YoEX9OsCuoY7mZeE+pyvTJJQK
0USgE4BtsvBXuqMJgPkSD52TiGRC/qMPlajByyWnWT1O48wMxLkZL/f11iMiYh/s
jDXCRpGY2SlpDbuoz/syGrQhJa8j8Em0UR1ROsN+MycQp3Itc771T0VPkfCpqQ6y
4Ns32AIzLaIMbnujD6xrNM56sp2rsbYmhG57BBUArx6dllEGQnrj74QaPplGzS4/
ghz4k6c9qDpRCy8vLkaSgunbOrTayfSZa40+bcUmeaE72OKZ77ApzJmFun8r2cfG
kIlScaV4cLr9lMKMrjQjVm+MYDFzDDH8BW5NWMKTjhiHkZB+wDXx0drH3SPp++8l
SrS3kLAwHippimY7GY4/gQk8ttimWD5yEFg5gQ0ZfCRwX3NGC+fqTbNkXk4PqXbq
NrfxH7GpgyBNut7KndIeFksun43m4S4RKdJLI59ve2YQ2/SjCfydnDn7UTMh9045
s9UGskpTMkwcpSZqMbzZke1mpfQYRJpZsyLIa00+bpyoZcVReEhL+j4uNNP1gPmf
rN/OFzc+YoqB7Y/VsT+OHCvE8CWlkqc470N6av5v3Y+dYEEx+14JT1aivSmarmo/
84rludyjYvJpyhyDUJ6S8hXFCNKUpHueDpFIqN2px+IZo/s7AfA76iDVCJNlSe7o
E3S584ucizMdRBNAd78PojxbkEpqHtVV2djxqutqHDxqUFkMG7JW0iyTCuaz06vF
iRVq+qlbwq2fJWTnVJBGzjcOkxusRn41xnVSmRzRNHo1RV1AIJfFZ7rYd8WyVOcg
EWptycF4xfwp30cxEUwF5kwr7efJ7QCLXpJt2qfP7lq323kxYBVgn4dMaYdcKosE
aMGljl/WzkusyEThMWARvEwAyyyp8siWiJn0XOesbsYh7NU+tvr8UrMYGINfkfRo
2F09eYCN2ocZGLH4xxZzo7DMn+sP3f4el5P+fDhrvvPrI03qbRGK401i94MCc3m/
PJiYWO5guzCsyNvU7qO0XtNacuH6l8fIsNjK1f2gaS0xnj6tHxJI9Htk8POAJJWp
e1uWWd3MA5g4b25Mz24mvCK0rYYEqJamudfGYL4dQQMIn/VjJNC4N2HpjgAldlvB
7brmaV0O/fLdr+PGbMsO02/xq0RYopmVD7ZdZa9Du6QavRYdqxnhxecVT6k8Rynr
BY5jaeYscdbgJTR3FAWpfS1o8dTMdGNINPrIuxDHTB8316CfTdNXuWwf8ZksTq2j
0QH9UYPnb7Fc1UG1Rt3fW2N5bbBHZAwQ4CXRd0gszTUAqrUpKk9NA8qBBjD+jw15
Pad861xpnNSZqpUrg4pUFzl5HUWOZwZG2w5lRxl0iZFoU8PG2dDiEdl8/1lxdIet
qKOWum4hftoLsx/+V+NfqExt6wYYQY7P38KTbzReK4kXnx3wLLvCnA0TiOpL6gLC
vMvYy0ghHSyIzYeuh7bNhsXs21+KcpW7KEJaUK50BbRPwJkU5Af0tNfegZ/AYKeN
pnWW9jaaw0OVMd2uv8BhmK8YCSAvVEUPit03TdAMBYmQMx0XJ2AL7lqO1QkAh6sE
8TN+TgSYJePmlfQojh7wjRZCfF7vFWNso5lsD5KDoUgkTiuLNTHBdxOVVwz1GkAr
v5QCGDiPbGN5qBsonLv+v/TjzCDn+/PlPK4q3WSjr82WlEeNMgksqlke6Fm2icZb
1FM83uRa2I9bfPUtv5DK3RV5u2XGBVjpEpj6NfcjORsSHUE3liRDLLRBemBtH8XE
BGsuxsqHsC/Xf9c+hnJtHJsFCMZjEzO52txyI5yd+CK+lwta/YppkL8PSuI7ULhd
qfdpDTHVs5wakzjxjsBOO1nqfcxEbSwhVEoCkt6BYkOc1cXSnqfbnDw924wxYngv
H0IHN1UgwEUXRo25qsxLbh/gs6FKEU8wp+98WCVnjp/bi+rvnQp3Od7bRSV2tU1s
W7I5DeTaOYfgDfagQwEZUqDA8b5UMh1WNQl3yhpljRXz4S6tgqbNGSqLSncI1sPR
9ateWbwc2pbI3Vhcs6Vp8kagIJ8KMWPGOhSJlQbweEfG/48fhoRr/0DNvWBAoV8t
xWq780zWeE8/AeKR1oxsjsWh2YxvLrVeZYRAKCbDaqNiD6Bod8QBcmeUCWWA+OMs
zW1MOPO3YGvqsXv9fcM2fKaXnF3gdHQCKJPXWrZhX3pItXNRS0fT59v77cPoctsU
i773PHYHvi0LdmC6qA2Tn3fhLEUsg4c3hIYK1rSYJFEvjD6dT6EDi5sdruITBIVv
kQliJXOYAJWFRkubrR973jRpDjzFIhJKEEQcPVd5Zvz/ACQvxQghifIP9vB5uq+t
2zpyMYJYTj1MYh5dh7QshgT/Jv0U7FhVPuyCTpa3ZkG6k4MSX4Y0bXnVCqxUFvbL
d9duPSIDToohnS7y45i831GR5bRtqaQV01HDy/qCWErGutxam18VVWWYQa9uRgBi
lbdOPLKbifojiVsgDHTlW5L4fD0M5HImq6NHD1Bv3r1p5aQ7TdAhdOgjaA/Ndee5
ythUNlLXRL0x2wUsDKJnhvIlDhEAqQ4Tj6L8AslP/5zqUptoiuSwHscrzv+Q8ymZ
S3QC+7E/OPJz0hzMYqTSjmzvwbE9EAgSpWmP2MSaLrAgY43XGLE4LM1ZpU0xTcM1
1g07GbTwFG22l9lgFox/cvCR+0fWToUIIaSmN87nW8vw7iGOy17NMzaDFOcp+32y
8JJhneFb4jKteNzdKK4n2ASqtU1DAYy2Eg50ylHveBE0nWWieMSzSG1C4/tArX1M
Nlocse6JwlxZuicJ21oCNQ5lEsBNFLt6AJqnTpKTgvBIsDIwHVVK4J4mSJIQbQq6
Tp5o0dflKwSyS6bvP5CiJ3Eb/TxPQk3P8jlHMyR0OAQIbmYmX3LgtYOLKdCuFq1r
zIn4/rd6MqfVrhdkl3Zs/DVE/5AO7WmDCgM4o0P0mDwiuPbYgihRjWr9KQvz3rLB
swWfspoNBI+BGugn4h5Dbn6ie0OPU5b8AaVqxaBDcHfn/fp80A9pVq/dTSuPvfXE
ultmDerOigq1GDw4yWR4D/W9C7ttxzeQjy58NwTSYsHqh44Ot3NHhNa8ZIuIMop1
L4wM2xx7vRcSjm1qpez8cg==
`pragma protect end_protected
