// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:49 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Xu4tOzCYfyeD96Bg1ifPD/C7CklsMKXvkrv4gCqxHhuMbgAx3izu/csR2LP1X8x0
jGizceup29GYAWPHatAecT5271glSds8flTietGq5xw/ly9hu6z5jRyCPzhPtsuK
S6PO5FV6rGwDJf15hHRAWNaQhrbA++AofSAYH/hnik0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11728)
DGclZAPVkRGlpg99l87e30wTCjNnnwp50b9MQG2zZwWodL7hT64mJ2FZQbQeaMHq
nvNgcaQ2Wj4mzeg1sVEGeYj28adkAoM44mPCRF5sgU7NQJVva0tkr31W/QZbgChc
8wscJPqBwr3qNomWBtK0gGWtvRrWfXXhBW4HlzPce7d/tYkts2x2BfEz4+YzB+G6
PnaiHuB1eI5hfA2tPSrjypcsfjvOGVhhDEBselsOaMaV1h4RwU5lhUSIxLBWRm6l
zhTCeN9poRlRWjwFggW/FABtC904GiS0G1r6dsxORdfSDMIr+MvVSqkMYYXtD2/F
JHdKXNqN6r9GfKl2fU8qiJzGxX8R2+eAeekxAQwHECxix11tqbTROlXU1HdzzHoA
FPfmN4NBUoBfchH7zjp6dTHRSF+VTrIzHARD3m6FqOXl/OrHcl5wipqhiMHv3uzD
MkhgQ8bd8tAfb+9Fc4tJxUgKIrtXkGlUJwZR1SI6MpasWijtnto759DkFjqRaDmL
C4FpHIU6ECR4JqmsuheytwW5NdmW+o/I4EXCR5iDO2qohU7pXAn0q5Di12TmNJVk
VulKJCvwtidinabCxuHER+EgrSZw6IB1PoT0fLOm/31UWFbwqBHQZOx+ldTP1u1m
Wa4/XUl5A9gmNuNqet3lOIewsY4jmzjHrYF9fh3WHi4etoALAtBmm3Ns5v9O89RM
jDe04SLs2gAoLnSxanLCxTrWhC2ngiXf+vodCXBO6FjQhejNqgCXh2sIpl1SSXdn
GEpzNZ3qQ9vxwdkFSQ/8CdnhoN0qp0foMRJwNvbBWd3MTxXEQT0wM5GIXQDmz8Hn
+tIqFFfE4nHuSG/L7nj3+sqSOaA/ooIPwKYGp28Hi2kaMODU3ML5l4BY+cRTIoNK
va2yXqZ2M/mQCgO0qwd/Vt9RFpx1oIY+0TBsrJXJcCcVGShR3BFNtGtmhfe5+Tzu
VdXJHAXR7zXaFMKbg6gmceVyFZcbcAHqV17n5Xey+RJqIIfZ1bPb+yQpRp9jfyO0
PHgcGjBmhOM8XRaPhiI8kBlR6djzZ2CQBSKaZggAzMJymPy2xC4SHIBBWfB7jsUG
ijsKd74egprSHj0s9FGa9mvpUx33T2uC3lMEiJ983oI1U3SYKW64+kExRB62xjUh
CT55FLXuJtL8ijEkDrovC5OE+oNcEfiHNyLXhWoQeMV2ANVBsc/rsA6tVn0MtTL0
w2ZpnezXm3YKMYoBTFk+nC66jCuxNmy3AgFMUMll/hY+CMD5uFcJqJB30YiUC4Qc
zUk8v1rFNvhE0OOt29mnO2vRiVzNkD638hrdn9RujF7BfBAhaOqGs/UswAB6m/sa
h9/j/s2U16YSvJ9Zq2UBqP8DXhEi4TEoSclzTjcEKOt3KYCwB/SR6zpqcSWkGw8S
EegqyfWAbyvSDlZ9IW8QQVjNCdyossqMDOK+BuSRwZfZgcwS2mD4P4McqOT4l6T3
46Soo661NtWZoXFIBzIxugkOsV+gJjLLzvVSIhe+xZRxkHJY9FJ5d+BUPosLfDwV
3d30jGu97ZTfsJrnl6ewTXhAnkBrmbMcv/4aHFepzfr4+gM1s3Mh39nxZiak+Pir
AUzlViywSrmSrEy7AHlf7SDuxE+dbx6A35ZVBJHxSbPpVwk/C9EYx1pN1Eena2Mm
BLrlUZpMU4nhTGUgzmT9+RJRrLdHvB9lw8d4GT01hrwux9khS/cEo9UeUMOUJ4Gr
TZLdXzQJ7KcsvKzWWPQgPPVcH5K8uLde/mEFbH5I5+9sFwfymwYK8/Zhxll4dZ2X
45N+kkVuoYWrI3sRR8HYtuTVmrD84lv3frw/qhhFTzobRD5kRe/kZb3c7tXZfJPQ
E5oW+E3z33Fd2bTeKRhpqCiYtDRycROUiNrZr6TLHgcLrl+6YZXvfacWJ6HkzO0V
EE+19p3YIjww0Vs4FGj+8D8c2DVoJZ9NSKGZfwp50lxjhOf4Ab7UIfc/VdIXQaOK
ugzPmNetIY2RsiMX+5OSIJZLEDnmhs0TmlcYirvycZYqWNt86Q5IdTuNJv/J5jwQ
b/rroI9NGm0s11t/0XAYgF6ehF6XZ6TXEIE+caE25YLYxVeRvQE9RtNx2VVr3Jpj
WuzFvp/tAWJCJuSF8KsGI3gQaKq27zN75qe11H6ER881/IDJP+EOLmfsY6GCPRvz
+c9H61Z09Vge32YEbNmG05pOie7sZ2gVg4mvLgsXbUiZfZoz2rPiSly/j19sTf2+
4qG2v/WYp3IYG7czip7xRO18nNr4rBSqmnJtgE2Tes6JAf3oyLdvePkdPY7LIrvT
wqdSaRySmiKxa0pC1J4usPwMfGmVEL5wRlkhNC1Ev/NAoStC2tdDfS++nVAX6e+D
50x27tq0MfLyZRdoNUmb+zmsWguY5sBe1T1PMMvcphP/W3zGMnIxIQoPB5fpAKtR
wb8Q53uLL6xDdaMbfzV9Ax8PYO01kkWX3lC7hG4vaxff7zAXHwd5NRhTq4V52Y5L
PS8pLmMsY/Tvhpx5RItgZ1XQf7gEa+np0jaspRtL/JhErMl09YpEPaWjTt3saqX7
a4B1R46nSdI34EPttHgrY3deFh78tM3HLXjjZ0X8vSwjm+gRNnWQ7o+XTodXq3PJ
s8+iqaGLybFg65jqaZRPv69R8DrExcmBr8emHZ3DrN4Bb7GrEXl5vii/Ajvs0D09
jk43VtoZVZWj3uj20c0w995TnXQn/5LQa7s8/BHMdx8p24sGJxSoBwVVIZC8jDOt
wxSOOvc3fP0GkbOdIFQ6xeQ4l54MTvEXvh5Bd7zj0VhMaNjBPjvPprTllJ+g58a2
79GYwl28IgybNCiCFwTIuR2f6f/WMQhrk4J/sOfsKCHiROmpBHXXE32IvaR9rzxN
Eel+cc8Nr4MgJsT3biA0DyM4X0ImCyXJjUoWVjMP+P9pjDPtykznHLh1oqiHrzK6
QpStjI00Eci2YoYRZMq14GPzj5vAjL4VNz+T0dAqZ1gecycBfG/PuhtyNU/hhQlV
kV1WiO2O44PlIJHHx51Cpmt+wW+1inHEmrJPJSKCZpCI1TzFuEmp0DgWYJf/fOiG
ERC3/Lr4JCnI9ypSIC202hhiLXbFUhfoIi4yF8MxKxDTF73IxyKcZ6sgJbX3HP++
Gg5DAdKFmUNwb3HetbaaMSPXFX/UhSPMj0Ug2Ct7xu1FyF+pDIXxwa1fQVm3cX5g
rcuqvrxcWTMbdEbfwAcbUAPAqu8Rmpi1dGkB69DpSODoxbPvJN6GgOurrYzbVfNW
CDEp/pAEp1gaFufE06Qipvag/8hiqZ42RBhdN/07pG7c679tIR8olkW6nfw1PjVI
86yc5FVgX1NKLHeo6Nlp5aQ/yGqiBn6HhzXMpm+XrIdfew+UXRE1UOyg6IIxyvKp
yNhasoCCQwpVseG3XR+VNBL/L7leYzoVmRve2jfsT+jT2kM+mmKLcPc4XdqTivHh
Q730tybahpIqJP9sbzyX+3n84+t9lgamlQAqvfFWLCsrJ7AjRVPup71au8cNB1QM
mSAo7t7w3Q4nm/UAEcJl6u7VERdwkM8geFfQ8XJ8uMRzd54VvOYvXaEet0BYauQf
rIOC1DR+qo1TeTPWozcrgfYdmqNxjsek4yiGOnT9R65DGvTRNEcJr+RsLJoqJiHV
POlUHN7hsq1mX6d6/4TMWLdvFbS2B7bIUK7BEX+rCExYNO2lRHy2sEoTAphC38Kp
HXUQ1MyJ8cprBX1rzUBKRuCCVcKz+hHGREUXu6X2eywUeD2gK2iz1PpElwAVXTc7
yoydtpeOdhuJPuosjlMgW92Gk/rv7o+fXxLIza2rfuzqAij69a9fJugUyIMFKLFv
8dkSEl42wj1SXKNssk6RfHNE5EL5u0PNyT671+akcOjs4F/wRvg/6lndfmrOOVdo
pWn8J5DvR0XwJRHfSatINpLGw7L3NkC73HPJNnIguTB61DJWefllajHhxIJw3xR+
KpTFoiQb8223eHvLHOS5aGeT4J+LhFVq9fRKeZFP4oDtGcJBD8eA0gZ01IWGEuvZ
Ac8un2A5BsEpac5INKXaTmd0XPxFCo11pMyYAvifmzITj4KvZ2kaer1ylalgojWh
qO57YRxkevaZkveL2vImZevpI+Lb4qBeW2uKDrBm64u4p8YdA/5t48eI6TRynk0V
31v6eop0TazUatH7+MpskV9irYXY1cY6p6sp19vh+bkJDJ/dKqc4MA6pjwfw+ODV
/rw7X3CzpGMqDOhtSTiphBnO/+3frXxSqZtxamNu9Bhyv5r/UDRvatFstX2QD4HU
2AicnfVJHgT5TzHJX49eBHF59kURFBVwMZzr9q5XBxMJvYr7P3sDPZVRhqvZuZeW
+oU8zCYWQb5Mn/7xzINRv+TMw0peI9wklogW+2XpABA7bMa7hdt+N6nPMWUumT2E
7RPHwCxi8dYGrwrzg5FzIhtYB/2QttbL5drpv1WYolR+AX1swmfDwT2PCdZfK23z
tqb7GO1hkhaclqDxNJDi0pYkrFOGpkcwgjS0wsK8JYgO9GMWNtvv/kLdvaXYMRts
ZzhZN6Rmusfz8rpVdZf4Z3RROKxyPZeCwqLAA2taOsLK2NhhDSzmN0UoMrrD/AMY
vCJOvi+HsV+CFzWxQgjXuI92rKo7j2LAEm9M/dTewLUiYiMZdJahxRT0aNJtQbPR
M1eeU6aDS7cuzI944pfHo1UHbtLhahKKDtUPYQm6Xr/75MO61j7qrKWpFTxmQKXP
93KBck9luZD6T/GmAD24evlfVOwKQz9GoTXQEDfHSMDcWLlqLZhuxFgjoCjUKbF2
WBEHXqKi6Z8ftdnZw8Ps2LZ23+hLZD36qIwq07yuWWgn82UqyhgZ0riWCioTTmNe
f/fW+SBNPC3+fdc0FCCZ7Wl81DY3mbRyx/vgFDO2EslXatV5iQLp+bIXOvrdkuOx
m3GVu03h9emVy0pL64QM7nw7XI97R5zFZW+Rbt4gkcXrrMNtyucEE4RiOuAIWG38
dGXzPsskzgGy0VsNYBzquoUfr2032JfEBhwX8V0JQXP/IAmIV0ycFo/UTGMBSMCG
iNPhJ8/yS/7JdE72/+78Dtk7ccWw0SzcJ5h9ku6pr1Q70m8Cox0SOOhQESs/SpFD
CCwfmdPx+Tp8OHY7MWJYMjZ3z7dl45mRlOZcCw/kMX23Q/2ryS4CNkQRw6tt0Zx4
KryFs58pHlhqeloi/kqBWmYSCkYIrU5BzpSEU1LZ1ipgO/Kz+HQAELnGnLH/bXDt
XElp/rUCq9lvN8EYCzcxe5eRHI/ZYBke/tMvMjCMVtJUMG75M+GTdjhu+a0qd21C
jjeOH5K+x1o0HEmHlRcSNDuxymrX2/nCsCg+2bDHBR0IBUcYkAoJXRBo3wi5ueAD
fdemsrD8A9kLmm339ejT69F1P/pWvIW5/2z4EoHCwXgjyfk2IYwVRTlOpHHArFlT
MKhUFYy5wBbXNGu1Ep0D7wmQgfoFLQG+tG0v2jOT9vFsF5YwnWkhbcPv17clnYaW
CFz76yLs/UECDDq9846HJnJzgbN7n/IKD0ELzBh88Z2MYIG0yL25Ls6F3JD7k/i2
xJZ0om3pIxLkJcmK8Au6o+BuH8aGTAiIzAGgXQGHyBW9n4TyUQ5jB7P9BRPkla//
NOs8glRYOQatyng9DLCtWZvy8xjB0UtazcWUIQWXng5K7ArDmbEtUBo8KzQTCRQ3
uxd5jJvtC+5jXW6WVOL/SPOZQu3vWpy5Wuj+DgMDfd9NG01+dgXGAD4qcJxQ9to4
VeJiFJ4YwKKg3uCZYOx2aAAWarm77OWv4QdwEuraZ35Dx3om8JYTwHwHT6gQrVN1
U0GTh2aM/ahPEq8Zr77tOOyGm5X7xYc0DVgb1R8PeVbPJnkFnYg2wsZRrocrxvYQ
NMOoGDHp9xkMDTRrxvhly4/4EVq8MhNTu+205iOSLhKdANbQ5WdKrGkIN28kh1L7
eiTnu5Yrxs5EuWFHYm5Q5m9A00MSpf9wEJ0dn+QG07bCrp8js6LnxTo1yRY33+Na
WNeN+X1qkLTBvbtsvcyA1XqSV5uHLRV/8ZvxSD6mdsjz41wISXkJzvYjLeheLJfP
8sCn6S1mz5GGfOGG+lSxKy0V/qNbCB6oEqIvEBMuTq19OrpSf5orTuZulTxUI/3Z
fJHz6Qmhrsp27Y66B2IIN4Ms8FDtcqJ1Kb80w+Ps/6g843rlXGn0qNF08bXH9tvh
rrKr4M7xxcSPeo7gNzscR7+BL2CVfyMcb89hmct9ancnemThLUJz+ZejQ7NDcrdS
h/aqBEMORWr8CbZMSCTsJzgkx0tDROes6iz+v/ESGuxEg35UuY3s5uLQhdpbLzp3
4dWJeocV32r3o9qNPKwVgLBULIgQGwUbySckVjwRgCJG+ibp/thLU6vF1u0fbPrk
FAIHrP/zlB2jJPGeCDOqV7aEoLuwi6C1aPA6gNIEvV5cG/FkvgKnIcEFYH69M3Wi
oMFj2AYus1XRhxnge4fKo2S2hjO03aQ7zAzFQyMI4kJs59noykWOXZMCl+BtpGtL
eiFdzF21rb6RAgcH2jDQQw2PFqilNRYoB8778kY8ZuvhOG/Q1HOCWBRoi3PnUZf8
9ldbNhv9P+d468XzW13n5dHEwIrjNzDs0737hHMgmOFEQFPtASHxfT5XPQ/DMkAv
WkR6QpRxv/YdwkCwm+QhM6j5TJBd965xluXh/+qGS1Ii9PjhBhmerkRPfE6MgqiX
I9r/XFJnKlj3YsbmPkzfyGolRFl2k48BlhQQpLNCHJuygyM/Bw/5IH5Qt7VxtUlg
afZfmEWwO1e1Q3tUmziwOLD9Gh5/Zdu9jJWm257tVWtM8Tlv4R42MoZPohNEOLPd
MI76cjDjxMK59OG0f2m5HQKMJTG1trNpuE6RT6iuworqlR0m/hLWHUuVy6NP+5ZR
uVTGfIj/7coIeUsfTvgoDZ5NmNPpJ3pfHNQe3gl/z63gJPRhHZpTR2SxIMIT3ix2
9kV/fsdAhknmt4MbnSOyKU+uccQkDVu1DTWQuj9ambxpeqbsbvLgtv0HNgWCu7XW
8Xg6V/B/3ibRojFLD23nvFzsMQb5jam9wVhALcNsgC3LlpzzdR2P5VEEkm1wo0H3
IWl6ggXXEBP/lhLkD3PBA8D12TAHLcV2g59qAD5kfFY91VK9XNT5yVTqgQGsykaP
ijEf6pvXMVXKjGPEQwa9cvRLL892Q1UWWyu/Mahek5dsDhOK1/V9b3d1Uh7ZJn+7
k4QTw4DMyLOvf1zEnCxWRk3etcwipmOJRYtomCI5/HWDAUJ4qhY3Z3EyjIyBM0pj
ATPiscYjyXc2W/zqNu9oYk/fGtkQJ88eySZSQ6S27NhUiIXNtxSoi8srIJTxwta8
RcArRns/c31AzWtjnSqxCSsunY3mwe5Q+dDRszAWes+zW0FpJJCJZygDVjisg39U
D2AoKFSLsG5DW4ybFWtz0RlQm1Dbk81fqeRg7QPc77YAyMZGZMFMdczF71OuGcz2
dp2QWrQaXjs10zZIpMQ9TO5i76GjG43iI0tXKJ41YCaRuAn5iDFWp4L7DGa2Kqix
yuYwuqko3CpPxJXya/sxyjQobZMy1fqr2ScaSwIGlklmm2ZjjgY2jm+8aubOJ8J9
0r0b8Xx7YJtL/39/iC8wmdlXzaTw29rnvwb81tYPGqGJ82AJplG7VKPMFOQwX9IC
nSbaTv+d27SWYK++6fQivhOC+BVBgNQA5kH4vkQFKTft/UC6jKJ1yDPP0wT0PRVU
CGbRdCw7xgmdlsQgCThVkTc4Ntw4HBsRqVPGnpOByim7Rjd7KupoiDB04Z82CGYE
rt+rxLdktOp+HeKSCqxHNWgbFfc2E6fHUhhmEfln9HtWlLJTAV6VBVYS0ZbP0TzS
lwGMURNWwdctWQdeXloptvEWNH50ntZfuw7uqL9bP8vmhgYbPA/dvs4zEwHE/iB8
SGD+Rn02ZK3GvKLV79TYDvETE7pNyjJqJqEqzzM6La7wGE62V9YtgS1wZ3s6n0OE
/l4QZDDt5JDIpCRtY9WTZwPASO7y7KUEvfnVZ/a2wyGcKqW2YdvxMi3rJdaeJIW1
sQw52pet5P9YsWAhgnLxZYBdMGzVUBcOFXmg4TomczQbYpI1swC+U5x77ORLpC7z
L0EbCnuUJCQco3a3cFXsrWBSqD/B/B72KnVlV1xzYDD9lnQL14a4LCiDF8oMzQX8
4wmooPY7xXG5Yga1pP4DYgForV7+UZ3cqYGi/g17c7s7+rqT2tqB2u82sZNFwF8G
SUqH4jI+iDUIM2rj82SAAGHDel6PvBY2ujCOS95nCbWrOxVMrJr13s5LlLjj6zKj
BLHB9ZzR/nVHS6LApXh6eDkSH3pDETCSqOA7r2U17dQoYBx2xVdqUqLI1ngiU5fZ
8zMiip6e6RmsJlejdEEYJMAxk3S9JB5hmm3xlWEY/fefRIrXc9FdbjiH/2s3Zc/h
0iz1dz5efKI2uMQrWDmG4o+Mhv6ib/nao/T/zll0xSLxwrfSlKsscDIVcMSnaUtY
+W8KgIFlZ+7fuo+5ry/o9cNXwOiLy7uEYOEzUVKalcEaUgMaCYmiVYASIp4Vstqe
zfcwywJVR/5XYJR9rL/ydpU9m1d1RZG2+3YOjF8XYj0h2NyeLxcJ0nVN6SK9CYX1
QLDiVL6fVV5Hcu4XsnW5XajB3BoBuIHMNDTHWZmGGiAENG5C4EIgzrIM07Eh1Nta
jA6zN02GUf2xOaGr+MDJ5Shf5yotX2+Gc/+GJ9rGI98kd2pxTMkPkMgJtxXBXuv1
AYzZDr4zpGR77XQEGqcuCblZePcypnFQhVETKQ020qZUAkWW+D4wk5rTBxEh88/d
HXc7xh+R6FoKXYtc4Aie6HodIHfvXv4DI9ISNEYpF5R+YCoBr0x631xdMFT0TRCs
3Py0alzpKmDeowuf1GzvJJ/XjskbH9BpMO6nQ83L2gRRbDmnx7qyIAxZCBa8NifK
HCL0us1uJVpLnqvR0N66h0lOJQDfE3tjnLwn6YOX9LUjdQAaQ7MDRwJl9MZx+718
Hlxj6MyaEssaHwDbYL9p2/d+VMLGJeTqMWFxuf8xDnU2IwXjEry2Wfi/DNbMPYmr
OBd9Kpve9OIz9ZmJzfgLs/Abg4bs2OOgt/mbmFNbNFt/HpH5EzBCeHIolsxzYu9o
y2W3lFepWFjAHjFfpLP6CAAWspvzLMsXtJHIknf+lLcGi/XTMsixW6xSKb5C4rlZ
z0FXhUL7Gjj/ATQj5GzMQSDRQX5GXEd58WPBFQcnvFticTTHkW/+NldrdFCsQSOl
DFvPq+0Ea+WRNbbne8qbERg2APBnujlRLTZaV8Ayzfa94meo+ozRv9QDPF2BPpLo
mabTx/uN9+Sx8JtSHzNoiBdC/+6Sp/SH7OEcsd/kOSB+4ltxsNQg/eJqi4deAPN7
qnGP9YOoKc3fp80Q4LsM989qRdra14eX8D0GGF6JpjTu/Pe4esLl3l0H8rmciTkq
SlpLx8RdHoncaT65ac7RIepOyJwhrbTbqgD5KC7PPwBOMLZ3jNIoQU3pQf6zH2mc
mxqOY73q39a14qNF9vQQ9yh7+usj/NHZpP4IHNTvOn2XmRCfmL7siQZvJ17Pd85J
z1pHBW5sVcgvjfeCYxkEUdjyCsap7b6dohJuhdKtehTCdaXijgS3xgVJCN3o7yrK
fjCxlex5Fv1ujzIl5dlyzbzmcebhi9LBWpZJHbE7UJOUuz9BizGii6skzkzId9c1
owzETR+GJEPZ3EOoSnaGwMGvaCGT7XL7bhT6nT7Kt2tG2bLeVcp+f+/NTRe/RBxt
Xmsxf74tH4VEje6a8/n23FaHEzB7siHO2Iuo54jHNK7HaFa43WFXZNE7LMvowfDd
TTnfgB3J+fiu9uJCUMsKjGHwONegyxa3XuRQjdle+4c9wkWIO5g8Bn540c5LXWog
51eHYxDMOcfOu0CEE2fWA6MrP7a66IPgGcMpK3aUPQ6Bex/QG/OIwBvG4stbjLBk
vPfvPUefX3nXgAnhxl3HnSk++tej0SpWWERVayOFezbSUz9N7ZCOWo54b9j4llcm
OKm2a9FHTAna8MsiFjSUxHaNx4ViAg7CmxXOV/Jd8gAt5y+UjJbvralbE9VZMTIn
yyjghRHIUABdDWG0CeqNbK0Qs2jBb1PopBBLdT7Io6pjebm6HrgoBVxebCqc6FpS
0cRMjkiXDTeoxm1rtcU9j+tassrbAUXS+UW71Ol+Tq3Akb1gnRhof+Pty0EMsXNL
bKbGUqePpI2GzdwK4hAUxuV8gyDsFHNyIcFw0jefHTBI3oDZLI0p+64TyGQkYbcc
8YxZjsxTLSSnQdh6N1TPxJUp0493An9l3VMMSGWW16FTK3jPXfwQX1YaNuGX8Sqa
CMwo6j6J/MqUh2BDWuGiVkGRGBfexTwfUyUKGSpSKk7tIktf7qjHviwLdVN2HJ19
hSUPb1J0/azIcFURq4glOiOM2wqfc6zEspFjCMh1++3CvXaArYrt/C9F4zy98oW/
mrtS8rRZ+JBgIhqmKaco+NSWr1axVQS5u9HWP/IYaIgS8o3cG/H6zz6P+Y+PMAUa
u7o4rw9qt5vMOLgdYsALNZ923AnNRC1FnKFpFrhANL+UsQwv2JrhqeJz9hNC2GXc
tfCAVCtmjidQynP/be7rcKP+ex9bFG1DUynGkBXgDIEq4IcCLtAuG8wJdeNFkvSu
yVnxofy06f1HcBFIJSUAVcBq488qPXUBkW0v0zgRw721SHZYBUIOHciAIL6tj7g+
oInR1KphIMkP+cyRzI0CfrK8ijsupF5r33aJRAMGzt0uzy1uw9orxdqGFQi06sRv
BplxqUJkR5eUZ4aZDnNeKWYsS1eY4bwztW6SVF5VwFxashZ9bpNvy4muRr1rsZjR
pDKvZS2X3aQbTj/IcDQflDNbKeHTNupDbSpncanPM5pQQrVgsZ7tjnxGYMkmyvuZ
gg1d+bB9BZPxaOtW1p6FAxlTgNgV81nYjSGHfBVT6uTLO0Wymuf93lJo8EEIxJxU
4umtxU4FDd4xtUfLdokQ7/oAhcJhyb4b4idgU5G4WB4UMr1BhAGd07TXPhLk4pHp
/B+rtHK+j5HNk+2ez6iUEHYkZpgOKXN3GXWgRdsPTe1Zr54UtyGNYFZAWyjIG1YE
kV9h3bqa69jQddUtAhrLAogCUqxdhfy+FZtSERjidzUiMQmsbEk5I7DoiEPwtonO
DjVg13v4jzRBxniXucGc68bptmrLurmM/wx+13heGSnQEvMyfDqwzk1HICv8wxmx
HYjbZxiXjR2zL8ThcmDl2Ap1lXKTJuBQzI/ZOcSnnfL65d8uVSrAsIYvIC4lcCFz
WpIWCiuuMlTwIdSyriiWM3I2L4W3l71JHvbMb9vh3GthRqLZH94oBj1rJYes2UmB
8ywBvkCQfFIBirZSLYBMHTxztvGiRfQcqTORKkfaVBPWX1k1HaQdTu1+M+Ksfyt8
AM80QK+GSXd7O+NbLXo97Y7qozoNp1rBFIaDrG8fUcTFdwctmbYoyf71h0FtV+dQ
Om2fQzVP1OGUY/B8aPJgQh1rFCHHIPMAa5e5+5RlsDSIRl3Nm1vscYRtcANqhNnJ
uhdtA7YwC8b05RbArfKxmY+CJJ6TTAidft6dFDLCvHKwlOw0ziW/q0GaFlSlr1r/
9kzpR0Eyl5Y4Fx3QYBr2IE9ljM6xpzKZfuc2SSG3c3kx2BBDQg+1w7LdFiaN3CXm
O4CkRy4J88B6eeHDMaHZYOI3bUF/qADHmWm4WBuPlqOX150Rm12+yGD6k5XHXECP
zm13aVxzSXTJVmLbEoMMXxn1afTsgZ42MdyRJLTZumn/736y9fBclGpg1JZ7rZ8x
sTx6O3OUHuGru0QrEtcHrdFRQmTto9nYgdquJHEa4r/LJ9hqwfsvXBoHBTF2VEMS
s3YOnIpvebcS/4T+eRBTCvXeRmJ7dRTzeCWjldXQTlqNsoyXkbbqZWF1aCqjNmCv
IVbDfDgd0BuYOoNoL0ywsjSC3zBofEHvhy7kztnn0HGTUfiXLQShgUB4s5HZTxgq
6DQqjHdozUWQlW4wEE4NvVMSH8x/l++FZvhyMaI3OPn+8jSygOJqCJsYoRUS+1A5
6PJWDWiPYJCXe97K43nOrToUw95hSlbG18/94EOWW0AYX7PPgXOTkwYPv3UVxXfd
OWVJGuu0FUWRw3NFyeqgmYm3eA7LsKE2Hs+fmHlxULYt2jr+xYf25N4Tm88vp+h1
TsOJ3LDqV0QKsONj0LK/K+95Ko1/lbuIFEbhnF2d+cX1XCKHQLuSeZxKmqoHV+HH
5cvjTItkNQrHWmZHay8DAxR/K5K1rbEhmxgh0Wrr3rumDmV8HkJEb7RUoTkradF7
+78he+yutITZWn/t9GFwhCoDTKX1u9Jb7LaizkKIkX0apcpV1mp8leWa4Z24Z9Ye
xICHbDE2qQBumuVYiLCIwaGRJrpCQXtmOaG6EzT2NEd6mSipgsMd9jKje7j36ZW6
ojT6LLWaXdAuieKcXoQOYW1ni8BL6XUUMdXDvMB0gz2YStaAf6PLwmoi5O8nbEuV
wws6yP6ApCCjWl6TiZuudZ8EYqOK+kuL+IG2rmM4WQp4ltQOMWN3kxQMvaORLyGY
J9+A90GbFDqNtghTddPrkrrxnOA9ZneJUXbmmYsTiWjIWyLtNcseDNn7i2pdlaAh
pmBICc5XSQ/fnOXsvACbu/8zgisL+F3BncaPS9ppjGv+xveC54r0o6oLVfMLIq4b
J1XEzVsEyIDBm2dDTQHk5NvkvsarDpjeLnizNAN8oTZormEcZ1I39K3SiGhoJNDz
gBGtJrLPDPHDKUpht7nb4mHMHErsSS6yd1uv27oYOId+BM2WvtLypxeRU61Onyh9
u8QehApJbLamX/BiSh1WZaqcdbM5gpSLYxvvJ1V8EdM44D9Dz3gknZnWBG4WyCXU
EMtbBNHFdJ/dcK/ON1swmiMVn4OejUSWfmzaQXlwtKL9u4R1TuRtC+8eBa6PB47E
wZZX3T2klZETs5gVMPQ6TPVTJtLv0ZEAFnTF2mGWUvdS7TiKBpqvDNXCLj+AGM+1
UODjr7MNknAQ4Yg4iS4gM/mAON0bEf07WH3NMnCIlWKujC2DSa6vfpXADT9ZZwgZ
4DgRJ1GGl8/amQqYbzrwh5OGFUETHjdELIZ3Tn3aAk+HP6rDbvzainUnEZ+pRZwd
emOHIEcL/BbuDJcKlT1BdOD64l5gpw6AkkcnUGRrAO3RPptKlm6C7kuZy9pIGd7W
4i4vGZ5IDzCuljmOBhbLTKDZa3lpE+dNxeo47QZX9Wuds4maimvG4dnr5r8s4hmE
lfoTHFvj25jwhYHbyRwQNkcJLV1jyorhVidqPd+xfmPgV0d9AbayQ9T73L39E06F
nBZNrpigK9AtFlAFM43rheoQN0hsH/JN7cXonE8l4orhGAHjCmREP1Itof2Fj93w
H2CSEGlQjBVdcKhIRoTaMw/Vi6cO3jei+uv6TSI1A2Sa3t8iJ0tAe+48eGqB1K16
UrGKS3JnkqlQkLCbjKLECa1hIDlrxnP2aMqMnMtd9bu1a8jzHBNNF5csvkAqe6zp
AXp9t2x0FrVv9gapwyrjR1NqVJZkZvQY0mxbUnTXscCw8hNyR1cKcSeqZHNKfHIz
fdcQRELzJ28MdwDXe1vvD7OUa27+4IQQjaHP5/VCgSjPwfgOkEUuPDI7fxR5+87Z
w03/Sfsnnr5iFlh2bvPhB8RR3Lj+fsLv7EH0/d+0JXUl1r/iKygSaH2R0jCKg2Ye
Lo3hG56vJyziBf/hBir7jg5J9EFsE8Sh1vsLtQIWIXWMI9mXEa3WQIMusMX/5+oR
4WB/0fVZuvpMacdkehN4di/94lROOIxZkzCRiL0Ng20nNU/bWO5Y2HMSKYfqBzff
XIyAlpSc3DZ72sxbhpGWvyahWPqnNw08H3y/gGr2KAjxIp7pMyJutIcGuyMf1aLt
LD4kIT1k+Mz29lWIv46pUBBLhZfNnw1UWMrHXon4rgZI3ZAW4mLzw5w+NApAB6+x
xwd+DVO9R1x+ArC05r40e0C+E00u+iPqLidTSoJv3EgmHwDgicWuFqH/5QzhI4+S
i1yq6v7Kt9RtRvLRCNldW/LuuFpAnNZ1bd6lTkgSZJWMQk3QXIexHXonqKCcOxwF
Kn/EtUnhKs3QTUokbZd6KgnRL612AlcnAJ6VuPuxB6yULAlt3ASvZu4g+TN6TO2K
r9RYK7cfPeDBUgUM6qybzdNvWKELQKi/Mf2jkQH1lpp8OZweGNmmZJ6682iGjrKg
pVzKSWkPUaKdX97JbUkVDylWuU9vAXx5cyxBlliQB6QDdf9NczycKfXBcfxx31b0
RN6Iw7kH0ZywDurQTIMIItVJlvKzyvaKX27dWel7xF1mLNRQI/Dvh9LeoVFxWxWZ
zZmkBD1GxnFS1dDX9lCm2EVRUxK9CiJ8zFyBN5dbH05xMpQPz1RMrT8XnMIJjiEh
3S9bY8DaeH2/MEKyRQslc2mJBxKnHgSwk4CAeq1Veh6eEH7VpcwzPlAvdT6539b/
6ReAjhFafRnWMawWxauHb9TQQrcsoGpmDBRZFUHC18XJ2+Ko1gxxUl4+fjb0I7eX
mhrUZQUBWyXBVaxHhOHmVhZoYqMjtdvxn/ln/wdHrBcXN7RWQVvwt3Ebg/WQNiJ+
xBJJDhqPByF5JyHkIgiJGQ8acFRrxzaK4kAUZAyCIAHjl7EcixcE1tbcTvA06zpI
H2t+NYApyPE1arhRSN+YWeawhC8vog3xNWvMGNuQcViTy5+eWbsg9CqBn5Q+yeuI
d6xY2xxHAh1XjHkTAbWZXTTV11S8xQTrQ8j92pI/YlH8FkUlPTR9rEw5FOnxHlAG
ywFIh3FAGbiG2y8nI8ec7Pf3JqK0MHLVCAA9qs+/36sIZKhgqwJcX8wmiANnwZQc
fSHEBP7YAgU+MO6i0A19V11lCGgg5CkPp1+78CC2ySDtoU8TivIOhCTTStLvH/k7
b8YTa7qaeX/NIuK60zo7hnDRlKaHvwEfvcnAuXAdmyktjQ9ab/Ptt68v7s5VAUsQ
JEnDN8fLM4hJEelWafoPG5EwKuZGe98nx9tYYMLL3CMcXFIPJgB3PmgGFW/womWj
gXqX3hJ/2r5ktGhAK5scIP847EQqJhGL/ym7EXS6a6AZ4e0wXiLxBt09TMbJ/LCh
vgZdFdR2P3qFPMleqWOGR31WeRuUML3tG94hGAEKiSU82TFq1BP+txKRwXwG9pOV
kSFhiqM2S5e8gtHxo3rLGaaNH8xCVEqA7+QHbvneU49QdF4UbDAxkcbUyTBIo76T
+eyFh+NV8uFGveKc6o5VLOCSyRmEvL7Bj9PTP/kQnGgBpuPmT/e3feKO1DGbDWPn
07w0ofj3FHF3B0FfAPjp395sDsZ81r4E2YcZnS0ikx90O35+E6Ebc95LjoIzq+Mh
iGZEfTFqeoA/nBgCcMyWRJAfFZoksCgFbe6V7IOJNo4KERY5F8Un+UdtimnEajHM
OoTxqWsNVkGzwBGGmzxHipC5gITe8//OK+L8YqrGEMLpy3pypqiPy/HZnohvhUVL
3nn6YPbUB83pG1yO1v+V2JWyMPhFALCPzkVt5FBWAgXgW+Z7Zw4QxmsSSR2RTC3i
mJ3B/G7BGZxmuHNNzD0a+g==
`pragma protect end_protected
