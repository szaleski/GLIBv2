// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:49 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
LzD1COh7HncduK33BPH79DuimFci8gTOE84hK+WDsXmDWPnltHMbFqlS4l97gGVd
iDwCPebtkkJQXZ7TCDKp94bYgAI8jyVFKJBAQWQufSaw80Rsy5gZ9SZ2hQ7OJhjZ
cZ2Do9XPmHjESQDfiV5eB57Sd15OD411x+DJinrWfBg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 2416)
ZNEZq16iQuU5PMUvKP9M/uVJpEXRpF6yleYhjdA24QbwEG/HeMAESZGrPp/TaNMh
GKQn04OCy1ZPjcHRhD6Rp/AWAA3Xbib5Kn2tuC5f4GjSPoBNtgwe6Zt2ppexNK+N
Hm9InbTE5oD6pQ7vwI4vr/j4VWytyM7/BflUbSw2SWfSAn9aI/nmq1Gu55FCdAeF
o88vgRLHsHmsN4+CcBz6LaB+luz+fEUeovuOus6rStuy6Fn+6ZjLHqCgGH8tDwjM
UV5ZELsRdYF0hjFlcd6Mj1B5nU+y+5tIZA/3lGO76TUNO9k0ULRuJ+7GIkUNAbaJ
jSoRk55P52Th+kVSDVlQH/eeY5vcycytt4KeEfEeqzpd2uv1MjIAiGds1T7pVJar
gjIUtsHabucCkQ7tOYPYJUzaVScAcftzWKmjzS9A7ZUnEGmGruaWU63D/nCLGmPi
VHyMQ5QVpGkjxacvfprqiJvm/AmXeg9KqzgfIclgi19CLaYMW1YOJJgdekK7ybAF
HHH5LHNd3AAvHCqE7Z5vwqp/2FDUb56VGF80H17dGURjfQilgqdRjwl8EIlaodyy
IM/HONWIT7fDZnmtuj/pmfdHnWaXSkCEAnclBXv/Bi20uaw2WmxFzF/t+O/KOzRu
36gkdUMCxjKAkEeYhQFtmZm4Atm1ar9rVh22t0cbC1u/9K1HsEIjAk5HaNiVYG+T
wOczkne6GG3/JzeZ3vk23LF3DjwOXepCqEApBUyQeyr5Px8Hpti2kd4ouFJ5atxT
HeE6YvnWr7q5RNdNaqvHEeqCbl3xwxNnYrcHyjjp9oUOqnBFxZ7PUWxT4jXfEJzT
BVcRz2yPv/Se+/idyT5jfUKy/PX2jLOk0rkku6Hhi1vjzskyu1Z3XStOgysUjGBv
YFhNg7Gp9f2v1EqERtzEtg6XqwlO+kHS+tNbjQMheUH53sB685SkTUBqbfzltL0J
EFvyHfU8ClDmrD3d7St2z2OqkWuPf2scxKva2l0+Ae/a8zLBRsTZz+PXLxXaqgCW
O3WMcrYMC9LJROnCwRTwdz05xNbXwJVv9QNRpPBE3EnQgvLWLgfpEax0OSGoLuI7
Dq4DnqGJqHkfjDNj4iTaNFi4NLEkJHYarHaxMneao/Ab+kEY94/fDZRqAvZ39vq7
aglR5NvUzbgxCqZZFXbnQTN5/AsSuuiOVElLADGxIvbTfDitHhhaMhJOOsevVSAS
o8x7Lid6x1ZY4B0AZI0NrvWaaoa0bBNXyRc/8k948vpHl9wKuP5FDQ+KQFmnoFCh
a/Ybq/FvMyjf8k4h2uOgqLs/FXBEElwRhIYSdnPqwETmsw4FfUoK5ty/Y07J6Yuj
EwN0hA+K6hIbwzNEUJx9vG/3AdDg8hkYTzUwWQrtunoogZASqIde2Se1bIZ6gf13
9IjGgoTb6aa6vBcnt1uHuFuE0vlIkN0H88Tc57+Q7/k3Vt14Th1FhkN/ZiHaaUQl
Kx/gzHFyYoww/CbFV+0LJI7NvhNtBtFJJEpjzDpJBzoQ6mi7tS5XdXdOh107jKq9
ihLK5ISgJ4Z14syrLtZs72Ukl7DZPwnzeKthYdjyNUz7IGXLd1ZNr5D/n318L5yc
YKIDb0ZI97SEXYxEy5eDXgz9FETxoSryKbxy+IYGIpV+EoF5K00z4BMce5hpQUPH
sHm77A9TwpqCTwgdjpcCAKYCVHR4La65+rBq3a14kAkNsLYJtrFAEHp45vPq5LI8
SDiCyhX+aTSdmc/A+4ni/qCj2jGJSCYAezS0ttI3Sg/1hTjWskWaiPaT1DTqbp38
NUlnbI19KB+tMXHm/gT5tWqZfpv5yxQBCzW4GjrRoVlCSP4gO0lzTVxwCoqXMH87
Q0w+bWexDDTC1ETwXeTFccjkmsZJcId4NiXL9GhBmdhgK4F/q2l8Nskxrt3x1bWx
d1Ybz6YwfeWcanOm5Qr6KDbROsA/LXG4NNSmbEq3pAgi4gUf4R1yOYzHT1BJdnhn
P/WPmiXUp/toHOrftTGSoQ8WPp71NH5tXOJ/+htOkUYPU6O2RfdlWSIw9VsCtvPi
a4SBUWn6paXMdaeh0RpUTFx9P4aEton72gBeA20x2TfuJbYhmq0+lKZ3kQ9ewC/a
p3Xa3Fzzf3qxsvUVfX4+JtlIuOl+nH343lR/HTYqTh2I/OCzYV9L8ccUxFiHGahc
Tzv3doi8uexB/6+dXPdArsl7SrSaj0kZolpY3epDkvJ3jTlYY2KqGdf5mOgGnSpI
QbDV49+4CO2sD59NVFq6jobMcT6hMCBgCOTlwVIgxHmrzvBFs/Sr36LDxLORN/jT
EqYpeu5fO4nryvhEXQiA+oQ4Ky4e+Vksuwa+UaJ1SiFjnjSYk0NM6KbWFkQU2UbZ
rgkf/HoAEcuHIs5OcAMsZcF+bfMGoeFkILVhHO06jBEvC8unhTl7pPpHl3xlzla1
FgNjO1Qz4U8dwodbl4xlk6xBdzt08pqp82WbRo0ghUpUS4H03ySB/SMdoeFSLfu3
nHiRBDSWgsuCLBzF5JNggqDPD13BpsFwzFD6wzh4u3esvJJndDC8EsGLo2XkmuUt
xNRU+/a8AMR8I8SI3Rjw9CijEc6NiPJ4PiTscniXmlAyDqmOtutWr1C5bwnN31RE
/cDicz+CUz5C1ezNA9lVfC54qEWt3hZuZwhaWnKXy/oJqMSMWaYqhR06vVtjhawL
lyJ2Oy7nORmC/VpNnLzY9Ozk8DWDAQsKHhBgT52kIGGPjd9ziVVJfS7cKPQLtT6Q
Rd/BXuWCmUnhySURnGBu8Cn9dhswr3QP9Eh6UFVQQNWAGNJ1nNDhhAeEBMpwqf9y
pmyitBgQdHQ6iKVHYxmrJWeAHulSibYWJ1h/eHvCH4xaNCyMmd4Fc/EZBMJ9ralx
QuU2ouyEJ32GbZUe4Nx8ecBpUZDYxSFLMR7Q0We1xKhazVgZrHhDmS2Zb0+neVq3
f/ueOeeBy/u6A53Ua4tlrZB7QYd6aRZy8EA+PCwq07QOfcWFj+ivzWO1aVNP5mcg
z9wM0vp8ooHwcist9lV8gCA/TzrASCrU3MkeA3h7ls6C0s+R5fWtyy6eWScYO7xJ
6WC+W4Fbu9owED/oeASeSA5tDv2UCKKXrBIGtb/VkvC9sPyD6SvBAe05tLunT4cB
T2uuScD0sb3FQL9UkSIJnOjYUVdl94clzIN/rlWrBg8fuEkUT8Qslec4TH5xg6DY
YLMAqlFXXBaUIlyo2GbETw==
`pragma protect end_protected
