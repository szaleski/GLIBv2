// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:53 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
TMXj+gJLLoeynKdHOVOf3w0hcm+VLVz8M3SRlkO/agY9tBouSRVNo9PR64x1BRTU
+roJ8OPrtu58KS1H5dvfuMNldyZK2UNLc6qNBay9GRQGLBVG9TyrJ9JjatkXLIqF
OrWGAqvcqteQpMxlSw3Yr70h8iSwF0kxTfI/jT1iU3s=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 20496)
SgIyHE5ECsfs9PnhHLmtBMqmRMdsPKpDZE2Sn1hsz1S1vPrqdb3VQo+Z2/uwCarl
/kTLGAEbDHGzEfCzD6MPTsEgeyD5zfEp/96IxWpApXybPm/oZZDRVmO84+4Fhnf2
jF+ytNLAqa1v7PLk1E9gGkc80FRvoYgb2XhKsKbv0RAmWGalgn93WqypnmLP2K14
87Ffap7U31Bb+9zyJ1oD569bFeNv17uCuFh9MRab5V9VpNJLNBFZZp5g7y4dHXL/
k4gSAVOW3qvbor3+wLnaM1mQlWySM2L7AixkWATrnZJDcJ+xOjXxv+pAaRNsk2jT
68c2xgp0z6HiCXgcH9G3BwBVkNEhs3lPJXIvPA2h+JwAMVGpf/aYFwRnlw8vurRi
HKsjoWkl9JtUn7JS+iCNp1M4hxoqc9tkB5SYZBemntfgOMN/CucOoDSn+TAssIiN
yLNNJUKydqHdZ0oV6M1flf6Y6IClt1ZlUuqUeNWCcP2RFIgZWilcSmhMyOu8bHfv
rsrFcagUA6ZGjZvsb15NnTcz2hXyxx7aLUEgpwHEXXwsqRtLDnq+tfw0y3YIvs1j
fq2WnlXYKBArSwwH3kn9nmb6NIU6t3Q+d2ngYWIqrtAAyi/STsFONylqB6nMvAwR
bXSGQ8UaS9wc2dOeD5Zi2PHBf+XCOBKn/5p5wgIjzJBnGIztPURbEKDFXaTqcWQN
I7Z8r6Wu5qjtQ5MNmY26ikU9YsLIdcKancv6lA9w1+/14IVqQpyx0PdS+UMGlO3p
FZg15eDkgTYLUgLDzTOyfcXIWFlk/oGDQC89hbI9cyCBgPDtWMa+7jFOwEbCNznY
yE8e+Avsv/twgGokZu9ZEolTHVsDMLpzl4XtBFBVS5aoRqZgzbJfeEgV+soujsPJ
sVi0FISuCTNcrjgxy6hpVrAP1/MBLNisz9/OtmPQxOJyv5ZgR0E/XTslxDaKJeVT
B0rkD5hRI5tK4E1aquZ4uhhNRzyeSNrSIX9YJh5SwcAOHboKkojIi4ToMYhQUWqO
6nCJ9pRc0I5LiaEU3gfjaZfDjTgLZ+RivKrISbSthKl83qWYvIeExgDMdUtjrqen
WSvCdzwdhbok+l0UqrpyM1+ShMPoWGYP2n7sM7+zTHzV5bfYyVOSap5fWztyhJ01
Wr15/DmcyXj0ubmmlYi06o2RbQdpAItGdNmJRXq2QlHS78JfcWLgNn4/22i3d+bU
2gTq56ZuIS5cuwDXUZnKq58/giRP9Mq6oxRT7qoB9JXhlDPb5gFjAMxKOrZTRZXt
aTcrLesT3s475tXp3vQ5tkgvpHtirFeZp5H0VmU7xm3wuLnqG4Jllz6kADegPPVi
xY+ePKMMT+BjmGQafTYIUQGiEYaKtBUptgR+wPK7C2HQpr9srfVlYCVMloDiF6oL
33eFUTYJRl3XtXEM2YYmqUBLL0b530AAN2R7qJqU3+VUFp5ceMnsbckw3sNcJ0LC
TWof0ZzvTX+4Hsn015RQZ/WB/7oQqxRPMgu45fRQJGp9kbkrPvScgVRtuEDlgkcS
e1HLfTu8/pkq8mU4iH0ppSzNCjQpgbEQ5djo4m5RAtjCZnjTeuWYoF12nox1G9FE
NI0rCf/sPlzP6NyiuftjlMTfyTi6fsv/zsmiziX7lcbFiHBzHLflvOk7+B/hSsqK
6Y6IvX4joe7JzqPykfsND7WhotSy1zM/Ug61ietsBOsZUXgUkL+K4RJ82wjtT2x5
yJPxwyrY3psWWeb7eyzV3BUuwqB/UBwS6zr+AtgCdAFAQC2uptpiqhEY7Ckzh8EJ
LsT205LHgHDO9OTARc+nKTJBnVnsAI/JKZLWI/ewakB/7dPztlcgv40vFRDvPYx+
uLFpUmUdD3u1Ed+EH+D637mOnxGuJ91dUFn2clHbL3yxUJRR6gG+ssqcyR6oFhRM
V0/7VrQ9CmdTZKTCjyUYpNtZ8yUiOgK9AtxCkaqlcnhYjMPTaMvXqG7CPkLwzpJp
5hXbMop+4ZCRuD0MYTD+NnorAIvjtA5x5fMdsAfLmYyvJ1fH6IP+BwMff00NwPSZ
2VRhAbwPdRj22xjDaVEa7mW7n8uZwdKRGp5Yhm9+mFNT/p7yRpy+qFhgaxV67iK2
TkSJhXtzKUKVybEHqwrT18uuTP8azoCU19tb+kVR5L6hca8o18OXlBF2/l0sHI0R
xyUdSirEvxq2PVhK5bdnmqFGgmNPrJeUfjEV8MEyHqt51byTcdLVEJpg1hcoX7rh
+NMUA4qyAoemKICZqRZhK/5FTiMxTDyiAZPbKUjQh5zJ9JgezNPdIDow80iZiQyC
Yu37A72DtcZ5ODNiZ6NRXF8tfkS7IVWwnSnkxPfEVOTnv1JfweDqfvCavLbazUAx
SN2xwLblD81E1a9nkAFa4P6dszhUuhq0d3zeJ42dnZQeo2Nmmt6Hww/XHY5wJzrP
LajOmyf05mxFPn8IJOyqz9MxsY23LzqLWa1lQCgimpzggNuxKjQ1fPxG0Lx9LhiT
cqU2+qcHzX24BZQFj9qrGQxv3aioTYOL98ebI4kMJPSIr2MYMqiHi4AUT7GAU+TD
KnsJOKEn3nMTJwNTi5jcvvIINfsftya+S6PRoyFKxXA9upoY+RBOevARnCC/CRSV
9IPGjfHaXwH1+KaJoJIcj93D4ZjjCHvFjEyAzE7Ej11qdkAKsqjnPMzrLkzurpbB
UASZJmUjHGWLJOmSkC0hlpj/Z3k+cMu8FRba+CeNUm1rwAEq+P8nNiKMV9UOFgb+
m111Yd5xf/XY9wQ8OgKNt78ffwLk2z3cHURMjIVvUVuEDkMFc4sWK++5WwnwX3XG
U8CK9ktGAVtyXypOAdEhrgQ29g4b5hgVthfC43YEps38z1O1RofHue0CypGcLTKq
WTWkjHxzCBdrKqzHpqvljWF7CwMkdHhvPmiqvjAW5qdYfiM3LpZ45HmPSAxoY/tf
Rnvp1xM82TLcGGRfMvL1v+cne+A8dETLAvEA1HV/rMtRWvB4TaWz1B/IFZVcEwNu
CzgbyJeXPEmFyENqsh8GMzV30/n7N5L1FlDhro6bXDKJ09Rp3s0gxwoZZU4ZYRNl
LIqxlihK51dztNixgdJZ/1Gir2ZaNrySzTgYNuscSPpWN03cLB01AgMvxDh7PhBK
YdXx2YNyT9l9ceXcG704jBB+jlLC0BhbHM+kA7hincZQree0MBoNnD3MQfLlemOp
2dc1PPLO+da67QjU1/ibOH5R9ppTjQuabCgfyAYqfn+Z5orpvjDN1IXeo2uffXse
oll9nI29VLWx7gLX1obJoYem2cA2veGFZQnFInLKtV7t6CJDrDH0t97JzRc9AmxW
mmhO8O0gpfJN0tHgZpG4g3GPNZ4VB4WT1xONe/sEEZC56Y8O/3iMHwcju/yccLCl
u+KV8tVjT+jTcvl8ZAhfU0BtICxQvt2ETJA76xnyrBqD1ahqHuZb2WiL631Jiior
Romjfy8Nazq4AyBZCdkKoLDurPG7t7zeQTKFlw7Yn2/X3eWZacj25JiY3uQsk/dR
dLv5zEaG9Z8exI0xMO7OKi+XuLlvCXCiI2lCJ2hwPcV4JQooznc7E591EyRoPAeX
/6mkSefCEnw1CmEDuT2ZweQFanCHAuH/2bQ0lv+smjprQw596PuA9XoJcB1HA2Gw
aaLj8WR0aoXtxFtrp32xiEgHQrn3/vaETNpl5w16mxYuZJX3sL+7UO4HYKg4qb4q
YVUisD+Nsq/eMIo9MYH2BywyExMs4wc7/TLvZ8v61iW5xmSVR5MaxGpmGpEcqGNk
LmOAlJxfw/VJBdUylKJaxB5c0Ln2zgk42fMhQPpHsgW1wXM1yllaD+eM4EbjtlUs
TBDjozLzMKG1AKCcc6vUJKF2/VL2B2+Br/MmxyAx0YoRif3ebtFgT9JNOskf580A
NmM5267jVqf/s/4iLpQvji7QLvkExgBWGye7R5sr5xl8qIqVpCS0Ab9b0FWsxw4b
GCRn7A207xj59SwVeNU4PjBrYajPZcnvLr4y+vGVVJrY0fz2Yftar8Zy+p+9HdqM
lriVRpSeCOL2+HNjxMZte0SojmAi+zHHXvKT0EK3VhWDX9FBaEtt0wGUeemAooZW
4ASm200EqowKF86AD37ePsYesaX2TiXftS4iIRZuH5d9hfoCuwybcnR+2JQH6V12
8f3727EynzaNXykE3DUcAGGxHZvOIw3h9FzUBdBIOqh2lGNzSQL5ZJ4WKK/jmrhT
laNbE8YGs9u11fiu21lyJ6kEw8SIl5bgWLZTMKVR9gr3YV+DWhtMPPZOi0fJAqSA
k7Ut/vmr1JjWFlMxWsWRHRlADRxLd37ZwKqBtsZuQ799VyCheOgPun/MLj+qcBoy
Vhs92FeMdz9nt9S70F1l9yAZLXdnJY/Cn1r7sB1J6tnMVie2vfSF1XOxrqCtzgcP
VO8DDfzVrabobB0ZsyjrJtWFEWs93O+KreDoAyhy7HnpsT1fg6yKjToatQbWB/9u
L91dCdsskcI2QMvMJ8J/gCJMG+7L6JNTNyYbESQizzgSHTfaCa5QgZJij/bQ95QW
63lN49zlXWoOlQQB/8IxhzCstxL6Mc3l4IoRTiYWkxpMUuBM0snLOpNBEdbpUDp1
NkVCY6+6263QcE14zX+sVTZ8Ykq8v6oQsNuDUL18Y6qY0tY70MFBoPayQ283lpYl
fCYyJlSJBfZ4+ENuZH4Wzpo76bofsdgc2luiFhFyDXFzhSHe6tAWQb0WqXVq67lk
4dVjj9zO6yefs56WafDW8BvNdrCB/HQ4/qiH5JyBH9aRMJCzdJW99OYgjbSM7C2P
W+0MVzQUXfJNM/lBtHAtpp7RrVe0YUmTSE3Aw+72MhN3YqZJkC+T9ong/aOIEPsV
KOHd5EZ0ZACkaPDTrUxCUO5vtiSwSjSW0f9MOYyX79gQXKze8mxPlpk2jWh9weOm
6YLYcJ5hDMteESjIO1w1LC698ycW8nziqPWOkjhdKl8VHpqYhguere6tBLWmWAnb
BnrHIENk7sJwo86wdqmiAaN4YbDXAz83QbqgnMJ9wYd3CK4IxuKRToXgDic1xyCU
R6caSWYT8opZXCki3vSeUQr1DV1GqE4n8HLeGK9RiCPgdX08zupOakQrsNvxAChM
0jqNetUCsxtWJNtcPBWbFSMqxn2oW+TqqSSlUr3mgZ+guXVMGGNmzk/2F//zmaU3
7p+S9pkroruaUVE5t6P51MAqXTCPrdlfscThj6ECjs2IaRtKKoZ8ZzqAtMLfye2X
g1kUTJajrXWYPOTRu/+YZ05M8LO3OmpH+Z+GNkOzmD1vuzU0NTCUDYMUTa+QG1Tt
gO5mdPxOJnWBEQp+15Y5Y4taCktWt1XZ61N1qmHZTtc8odRFZLFSkBTr7+dj+ne7
V7y0VAtkiDgR1AIL4N0PvTXsJyIfPb0hMVoUY+9D40dw5M+HworqcHbv8QzsvPfH
bRsjUYAMyhZEPUYdplCM61jveuQGWlLwLKohgk19HtawXppBbhLW/Svb07tJImJh
IlhxhZw7cJNFkjwGokMN6I0HtZnntnDwHJ0u9alByCyZtaOJS2DIQ4Cuo7plhdLe
h85pnrfiR+3SFcJlDZVNBZJNfjL+5ioRgVNquBzWWo7VuC5qjI7k6ChC/ls5GTEQ
vpOeSHPoiUezC4huQKltBxiKkmt5uwhd9j33ZoVVmPh/GGoWKuK3jDX4v8Fakfoz
5hRNVNG7JZTHP4Vs/6+RLkjbvo1zvq/TzryU0jgs7TWb/5gOe7mo+Zko47qMZ4Ix
k28UChAXG2rWquV0AcImX2+TJC8zWqiWtlUFs5lBRj8w8lg9dC4f5sKRmMXkF0pd
sR+zQYP2kjmLrQk+fahfn/IVMwSrTBS5M82Q0af9DNBNSufPKS/T5IOUJgzX+Q2R
569+t1El6t/OiyOqfXe/GXO2VeUvAjv/3dFSCa0o6/EZu2P1mzPNoPqbNtOt+cKo
/mQvpNkHIkmXYP0REtf04gLfZG/V/aXFScrJVTzrnMQPREhs2SGMrRhtlOiUGKrV
szMYJA/QllVTH+fAKiXUtI9oA5suZ3rvWeHzgP/WS8/REe1xMxfDmOy7fp0EWLQU
xk33pl+I57brw/U3WEC+bh/kOjxGp8mkkL2RB56TQ1O7EAzwZtvqNunD5NztjP8A
81+cTJjzrQ8GISfoaC+mfLrnP6+hq9h74ETpEQwsD99XsDbWq4w1/PQ6aV9h2RiB
zk8BWAnxzNx7NfkelkAJmKf5Ns3qPpg6FlTEX5z4GGOauxHBxhPyCIlMZshhtq6l
v1vxx6M3wQ2lfI50Trm5+etBDKbZLzzM765QSVijApZVkODqsopcKbyADHRzuird
P7Vr+kFjwxxjck49TBfm7eUqZo2akPINRZ5FupEMJMKtneMQHDOHFYo8rnaH9ymJ
zTKOM3A/QDy+FFz6Iv3kdA3KiFyNgILqWNm09MczBuhwabk1XuvFtujdK8oq492y
MnpCDnG9aONulm1+47Z2yjJ0Hkh0PKIodmIGnWgV7SSXfNP4pWbCeuuY2Od0EDll
hirVM7ChuGI70aswWa3AS+H4akaKFF+/PYiOZbjJ8INcWhxU9smTgWVVfgYx3Jqz
E/gjnoelpZ8LZlrJG42PZOV6xx5vu83E3lVyCPwwBmd6QGUuOb21uIgpMGSzKySL
uMw0TpmySftIxAXwdEql+T+oaQ2B4Cr55OlSonN4hRvTH2SPdHNavfoYLJvAns1y
Jiu29iPqsqWfVk7JNwmjNgqhZgnuwcahOv92LVX0R3c/JlmYOqY+xs6OVhjNwPMQ
AxjpsoNLmv2rvq0Do7Ma2L0numhzCW1Z3UhiZa+mA5RX0BNEyo0Oub5JsODfIFi0
85D4HL/MrOTXv/LKcSYKa0CQ7dhvgp8XIwd547gSBiT45iKR7LqRtsPnA+9K1AC3
HHesYEt8jpnqYipBFnauDdDjTbz5KwnyeGTX/LqEuRqbgHNQGvfX14Tz3VMp31i7
qn6LXjbFhPTjxuT8AUaQ7QXkPy8xrqeYsw2mK6uDKQdRU5rA85VDt6WfFofOr/KX
D8jpv/WyJhzaNzJ2LdShDgfhwFJYqBERANKoGKaqqCTqe2ZGYJMGY1OVzic5qpkc
UJanZeLWinkiFoJwKzhawrrKJIFVXfk3R8K3R1iN0gSfFAanLIqBoanJhEWkjo+9
rBldk6EKDkrak+WVkmgXN1l+y/WJJwsT/p4qYV4oGHk+5h3Fu2Z3G7ELUd5r8QRu
CEjbt0NstwZYiAhnROGaAlgSgON6a23FBI+lYGyj7br7UnJHcmFZ+u4EDI0u9zgI
DuNYkKJ7arMsAckk/ajErWUO7puFXwyNI7CKZBJrbWXEfBqGffkMZoYOuE3RFLJY
KG7UXZSorwXjmUN+tywE6i/2JeJen9PmxvBNsyuEROahFRUhCQdI8YANESWP0+Ix
kz9LtJ2LI+/kfyFjWhsagmheULgERlDqvhH4DWeaOxBv/t2mC6DGPav/gm3Pi5kT
OiqDLpuHL46pXLJRaSNmdIi+t8RIuQ+2GqXSCF3sM7DSSmx6Eh+muSCRhOIyMiFW
8+fonrHXIhMJod2R/qBaTxQ/zK3ZMLVk7z8ti93ENs98hGLrNvu/kuBP37esyxao
Vc+CD7+43HVsW+COmU/k/0xGHVyQBsmIZ3l2kjQxCyVZDOD7uZILqdid9pXwkM4y
ftvAH7PwKQV+nnby5C2wRSx3U5I14/fd4PjAT97jJ/+nvJYIk0r5EaDLOnGglqIt
Bo62ihK+AK2IUmTNOwR40X0y93iE8p8RHzYC1iXfGb0/qIAQl0p9CpLdnmmLwDIA
rm5KlxLloqpZbJhQq2evbNd1NdQAYE8t1OIXnhgiOPitrFKKQDnPIzWnC5yIG8r9
7upBLOVhgPV7QsvDczfUz/e+cHT8RDFWKQ73ZivvGCvuO3o1up+hZFKoTB39txY+
pFTbzVF9jEixp7G6YjSr+xjEMhw7p4gyuYi6texbgTqMq29H/VezzvzzVMc12yec
6FoXKLx4olSI9mTBtr+i8T/TSRQqa4ej63miRR2odEDo1ZrUnFDN7LBxRAtVUcQe
NSjOk2uQUdtgLt7BqrNiGcSD14h17Tn/Y7USNyi/HQRVs668Rp2anfIN2B5jHgGk
IdCQdN5LK1wNlHD3xyeYlRELCYbdnbxt6IqS/a6GfN4KBoPhWUmG7PH2RPFGXKKk
C12e+A14JA+J3l8Alz9mm6h4gXucko1xLa5N/nb2Pm/kn8PNroBQXnXpkfxzeA2Q
IozCV/LSVtVNx93x83vDdLlVjzmBmq8q7hWs2h7T1xZa+88MsF1BDiaf4WNGC3CJ
YgQHl9JEfKwNjXKCpnNVN9oC3r6qdK43AYZsg2dvq5U3nH6qzElJ0fnHw85m3Y58
csrKNxSjQYfd5QibZZCyUg29uVU/UTepVVku2ly2DUOdOeTtYFkRdLrQrn7Fuh25
XHwxdUi8EfzYYkxifLSArbwjvdqzLppRGVGjcDtan4W6yTp3CUD3EFoKaXyznZ6E
qSEvONnjMIAfXf0bj6mEKbUGc6KYXrGU/+RKI9MItf2+PPrptno2AkTFYMbicFaW
+B+cl6aKnH24XqZwSjqGw5jnyHjoXPbx/qZUvH7+go5W1EqhZOAftTY1/o/5UXQ/
fVxU3E5bRQlsxYjA4Rekh3kmtZE/4PQhs+zvigGDPBkNimwOkyLwDmvWX8uK7X8t
UyLv3LoA6/WlfrmH9b2yA3xg4CCVdpbbyO7yIYwZOBLzmLj4uOP8XLWYVz4PQCPm
xvDnSRrIPUUHEMWlFLZo5Ngh360Bw63uHWozEYkEqrBj6CdxZWfRMFkFDVfk2Uj1
HCJdPmk1xjFs4ohoR82FyMCegveKxojg6sTZyF5tOIgXEG2PgjkNB/Zw6ZSFzhQu
3IsI0FLSrF4DoJ1B4SMijoKEZkL1wn4IRTF5xzDpMzVvPdVuIQTH+EueOTa5Prp+
SJurxxDcetQSvKbG6hmnTj0bCnTAYdsls91yT69BU/fJ9u3q1iQcvTX4bpDo2uOY
9jxWskZvroj/X7MwGxd6/kchlOEgE3WF8ZuJ1xHkP4arBx9bBeU/GpgT+7B736vc
daz98ZzRW5Q/jQZY7qRfvoksa1+7CbMkjlRI6MAKoBpOi76KMdHr2JI+Qk8MAHgb
BMbJVDUNmPYIMWHvr7Dqppd3X2L7o3Yhd5WpUIcAs4zsIPjKx1+FsSa11+Uhcmtj
nBbSwyqcse6qLDRoAFDV9kBXwtA1vF0SiBY8aGTaeuXypIv5Nn2B6JGUhhW203lP
l/d5XUqM8N+jyRgfEUQ0s4pjKToKF4VhbUo3WFOQezDFfDKq1DlBulz6t+5fk4n9
itNPggy3FfkUCIvmW52RapsenpwHRu7mbZdJqNm7ZfCg0EG0FAyQmYzh2QTFnicF
mAb5GILXozLdWDSjORhR6bKQ6Dfgbwx1gPYErfE0LqCJkQR3mehkpfgjBdvYJ5Cs
ewYRo7yqD9lEkZZ+D3PWIJLWlHWxEZjZHSmeYCYH190bvqLu0XIiaCLxEErpIoMi
248FdmORo80SJaK6B9LdnMmXbptQ7aLoV1aFN3R5q1/XS8VgKmYLljHY7jPETVLZ
IcWxXay5uFVH7jox+LXjIKBr8l2X5DPygGMb9DthN3Y4izkqVU1p2b4OCAKLcUM1
2xMQiE29bJlfV+mZiHILWud3q5zSQ/2Zns1n/e9Np4kTyHtAfEt7k6U3irDzLJbw
/BblwallQ56DKCAP1sHeClnaDkp829hIF6O3++6FA5cIW8nNcTKuMWSRM1WJpGYx
aSLysZRQH3vbWf9Y4HxMp7fHUhj0ClXVmeqMyK/eCb5bjQaTqNpQR0lMMsaU57J9
KSqwpIol1tpfaJbwXKojZhapy1yKazxqBaRj5VB4unGXZK3alWnYctl9FEhzJl+8
mUS/+6gUiQRlF0xui/G2+J8jAyEGEFlKS88w4/uppLx7Bwq6d8WeU3O29EpPKJBL
xOPh2yz1ZWzU978fs55XsRpRRi6Wan46lzenQt35Q8L0/LIho+1wK4ZQzjnqjMC5
Nb0MpFv3hFrnrfSGaP8RxjRIoWQ07ru/J+BkwtO6KwWV9gnkaYxjxC3zkgH3Wv23
tz0bKeOoqWz0Kl90aYozmNG5+3ZPriS80Vy7Cp6xw4FYtDNuUhq2hnH6gWWfC6nd
Y6kFYgNM4f2/QEaHl4yaEWtZ40PrXIbruwYKdBN/asmhEDC/n0Qfr2daZQJ6MDr7
5efeg9jWEZdyhFds4WGbotJEkH4yzOiS4T8an+JguAs+pj27ALYg/UxJWM5TvM8N
gkYU4OesOSIzdgBBr5e88oo0DW1e/FE8vaWNDvNnOsre85U0A0H8VKJeouwaCEHC
6hLXBgj15wSC4qlUKVZY8QBXYHxEVP6HloOZX500DP7PG+cSPud018oNpvUESbFd
6WLbVOLFPRqmsgfiYCMProy18C2uKnhtU0AK4VNvBbvXMEq8cB6mEji6ULeD3aFr
vdnxNR4Fk6cSAplyDNs6+GbQjJBab04mkxFYskMxuueSd6Te7bIE2q1Ai3aHR5cl
AYm4j38yv4RZREZmr8jh8CToltRomd7WS9ZOav6Zf1CD5cVtSl97aNPKKo9zXDre
9kOMpVCEDlAPVIVpMeeTfVQL1gRdPPiiIQ9wBfZQvQm0SPTLWFe3gDcErKiu6zus
4fFc8CJMqqu0uTnHNqEWjqQKpOP9svtP+Ksami8FQ2lZJZPqj6X7z4hdD7YKK2OI
lKg067uNw4X/WCZ3ok/s+fI/v2RcdX3TEPA4d5E9ataGkGfTz0yM2eJ9ZVuYxLhZ
Hg3UM8NWV4lH/p8Ko0P1B5X1dn/DfN6YPcm7tNpghgAK5ZN3mC+hdXjazrqmVHqZ
X3jnACEyEaLmfZfI72Mk+Qala7Dy9+PGimnsNZQSD3HiX/Xwi2WhXei8vTKWvl0t
Gdt6n9OKMR2Asn3jhD8/gUo+8SA84h48hL4jst4AMgaz71c/CcA5/BhCEfDmzGwx
7HDh/KjZKwB+AAvdixYU8ylAXYUC7/aJUiuQad7hq2GIRng87eUOXTU/BBs8Uvm7
tnjgZ4YXj4A6LJ+EUzK45uwJPmcbAiNkc+3ns4DiZcrh4wmx/0YTdUrHujJB2+Ox
dFndKGMZyzY1Kej4RZqI0Kwvz4qADV0j45rgchMQfEiyZ8cdHxlusef3NyO/ZXJ3
5H6ui8e1N4hELjClzoEjkTZG+YMliZSASjW9uOefFYFhmSSjJiTNn4878OJbedM2
7Gj34rb4UbJ4/J4e3xcljeFuimzhO2BFekiEw2szrSITOMMFpE5veZ110R3geLL0
l4HABx98Cck7nAUIIUWgItGE9C4z74BLOe6Yi6zppadNMNZ+FApuMV2mT/V6PHm4
7Z/yvVRnJF/H4cK058WUT0coEMItcIQcNRVdU/buPv2YNlVHoYvupWl/iyFyI31C
lsjo6iuTm9QUXeBmdKHE0PW64m2y9g9/lrm9KHC3zkDsW77X1374DwxRKxCm36pn
3kh/tzMvDgrDvvLeKGSA20oeiJUnw+EtHSYC9W8ZNYmbiMYYf9WMoNclsXtIXwkk
YFPEptF7LycP2I997a7C1chK1YLt+CRj8nYJ7FRWsOKfge3BE6BElmpJrMrjALKZ
WWBWfayRUau/fEaMMMLVxKs90RPalkOEMsk2/JhvjPl2i+qgJdpAZG0upQMSxmZD
DVRbC7UoeLtH/4zMNYiVzmS0ok1McZDjRNyI0ire/JB15bKrc9Qn1qgZ4MmK2Vfd
De3X1lKoMp8jsucLt0Asi7zhJVGl1shsw9oq+8Fr8V1hmXNcHT9E3EmyatpkES5y
Ua4uGVoRw07Ia++MJDu0A4GABFzQh6LgreaaR4UOKntmA/HHbIDI33eHUJQg5VCw
MoPdIAIPkynaDxfFWy+pkqb4JdEEK4YQ1UOjJM8uvl/jqpKiR0odzqM1maKxMqYJ
9F69XiTKaDVdNih1O5OoPo5hmBk0AL6aHZEeJegV8CZm3wjxnApxE1U+j+zlZVmx
+Wh+Sbv892UpjPC2rkJLBA4n+t1IwwzQr1j7PStS4R/rPDSfoarBkFE5mEoCkgBo
XJdk8FYfKMNCnuL4x4ZnHAqY11rIe6SMTNjTXBkn7QrdEWi72sSg0fMIvZTDhvQE
swZs6X9fihWt3j2sBNebLLbSF192NaP/LF8867iaTpT08rEGnVKGFGGfWaujl/fj
rauz+94zemqxug7lOzZC2IdZmmk9c1OgBrXb6GRXIGOWdsqybkVjY32WAEyijSTz
J25My0v3SBNkEB69VIOl9rVk8p09a++vrSVMThktf/7bqGw0ZVXREijVrwRrljnX
SU6kS29TxYkrO0wK06759INsM/V1PCWrSLQD8NTMWCHKk5DzqFyMJGBqE6jxOoHX
SgSt0difpO7wFfSH+mVDF62WG8ONyQKWmoE0Oyjz3WwrqK6TY3AGAO/RdMF3vOHj
rg8LaCOnmbLFQXVZ+WY4jLw82avVgebLZJUe0UgGJXDSl+NZ4Il/9YTTuUeLFcMP
NLe5cCfNqXKifTBn3B+cMmlJ8s6vc1kqJ/3dfO+LPEuLXvwe+4qOhzIxtE0SBbL9
RD45M1OUqAwdtJ17JJUhjNq0ztsMaAms+2nlqHiIBw8C59w2mtmT9eRs1jve+Lwd
lTfgdkFVx1amrQABnaQcLjP3RElulQOMv1yBTLxBUpMNZQSb/E+5bFHqkSBjBaeo
j4ylen3l/ljah7NiA4F1wRsAsWisZxzrfNs6TSvzwO9ZHWnX4AhdeQCC2uu5/9A0
VC7bnhKnPD5/Ut57Pge0RHRbeeeUQcLGE3GXACOYFNDbdBh7lWruVNTO6SV/Xxka
kNxc2polY3RTsEkNmap4ko4B+u7zodyo3BGPUx09QnrCk3WVP+as1lqYQwZFHhwu
WSUlDY9DP0NeOYiqTGBFEMS++LSGErFrudvAzZfowqCAQSVeqjb/SZNaBektyVTT
mRTx9QSayXXOuQeARpnE/SzNA/DmEzzpTPURdRo9JHWtb6UOwmpBeM/2WVs2BYUs
0TTtUnHDCXwzkC/uJpdsQBsPUQSLkysr8ecjwMrbUb9D9gTUa5byv8+K669gdxqi
p3Mvdbf/Uzxd+uTkEAW4TUPDOdEFmhMqiNUEL4XCfsYbiq//hKBxAQr4Va74uQCd
1+r34qJiwuACuR38l+jjSR5/Lgyyu9A74Z4K1uQhWIQEssSIuxgDUb9jrqGD29z+
kPegmY2QwnDoauFlJ/jysW4Sqo7kMGQ6/Q3JHGlmxBcr8FpOxbe7W/pT4juIiUdM
OzPuBlYbBxe6G53Ry1Vg951ruCgfYoQcQAJoLO7VBkWsiChu6r1nt0CrBX1cGkZi
bn8EWNQAF5mdQ+VpYnhfEus3niCfQ+1GxLOTEJmFGUirIPfRJArdM86c8niDYcTE
tNBAGdi5c8zFOyvqA68cA+LvTNACG3507YM8lkfT5H03et9ymZtwxJGm9bf2XRcu
b/w2pOoF6KOVlG3/8hrai5sG6PDxsOLFwb3/YBLyOKi/KR1jlC3c2AOSe0vPHn3N
DlFbURkh9unFsTq19MFm4o29pptAPGYo6wIBFZCXZSKd5rPcOmdeH8Q2tydEvfji
bavfmaugGH0/lVq9bRI1gQcJteYGz64ugBwURpBmLsKayy6NBNQSxXEew81Qb0ML
1QBCr0Ql/E7h1y9wML9rNqx/F/laMyTt6uoOmJniG2+48IDaf/OjDge0pWpLce6f
Ul09raxJX1L6J9qh6DBIE0zoVmRX10Z4dSqE4O8rXmsuk0hBTv9cWqRoxXOt2jAN
KI4dRagM0UJv4UYfOnYkTJmSE4DB0PrZOAz6+OtREffMZ9/ps9nUj0jNviWKmG7F
hYtniXzoerLKGVTFASsVqtDtvaT49IXyuRA2vmjwQMkHR2Xn77ixgvb/YsO3Ur9+
Le0f6BiDumaGDFllnn9DBQqfbeDOIkjO72ksfmz1k4E2/Nmeig7XyHvk5yXIJFIO
QIV+/BY6+d88qf8zjsZkZnzptDBp87Mnj04WVv+ywaW5+plILNT/xKnkfVzR60Pv
TO1OWz447s5U7oHTiIEU8Has6Bo/k2M7Ww1J+In1+LJqSHmR26sYERufLKzwRwmv
+ZjuCepD1kwaOW82tm4sNi68Py0SbLVoXtD4y/8jm/xR8ax6364cKyKTq+k7VJ56
jUXNpIy6YR9JaqHfjjrsrHh99GJdsZhVUraHy2YxLEoN7qXhyAsuOQk3YEJfpbJE
fLq98CNB2kDGi/n0DQ3xXi52n+uMFgt72ldSVqvbq8xDUBrT1qXnuS/AZmUyJMdc
kbQ8i7NG24XwxorHUKEPVBYkjNlZwWoRqOesaQqDf4j1NUVc8Rl7nQg3kVnJbZWQ
2YvBqiGssSkwdBPH440PeEWdW76NWXfaguB+EZnU3XNYkrRzmbs/1yEUlXZfl9n1
/x8dZQK/TPSah1CVQwf4hk3MpLftCukdeiJhY7NNdR52teNDPa3BLp741K2fqGs+
nB8X00GqBqVS7V9KtcOlwwqCEto20wwR9UR0n6YrfePp4FEOWs6+ZeERqxA/zukQ
ivjtVOHs7HInD95eLYivEwt/lvoPv6IYOWanl+XvPngLEFvqhTnWiqy3s9cioyhe
15FfDDUc54Qvg/R+qTnYDM1ZWEKoP+Bnb5xKEjvLRfB0JsQ++zMoFw1EIp4M3K//
YcQNJO1cjFP+KUiferzuHgNv6hNNJPyXvfJqFLYYZr4XAXS5a+iAimGkvrXSzx5w
p2Ln1xK90MQ22Hv5s10vznzkIfshqepDESsk28Tr5XQFAy/sKRPHHWk/QIF8H1h9
Q6w/ZHy47yzRbtY79soz/YLVY7NAa4DZpyIWlSQfyB9D1aQzw4C2kBsJ02jyNhqA
+mMuBb3hspYHx/cynqY+mdcx469kg2Y3P4+uhVwI1TTmlHSGyGcjkKa6c6InIZMN
rWhqrLHoN+Py6r9gjes3sva8Xxj8/3CV3ufoe8B37aCAQbuwZwCw1ofjL9qnH7zS
mBDgBPkcOBj212Oh0baQASC7Bs0UFvnalLtfpKTv9icPkx4w2tCa/Ex5gDWHMu/1
cB75awR550lsFPzUYiwhZXXeJN2OMEYePPKA1tJ+/IUrBBz6Ki/DQ8KOGAt1vtxi
iuHrdjnaFnWULJJc0hSNp+X52sFPwUlRIRU22bnmSmQ7pliaUrvJ0fFX2N3najCt
W6DIhAnwn2iCOi216J2TM9ZvLwNC/4SgeEkIf0YXCP1QIypiEV1ZxuTKxXiYe1mP
FIasQNcn9aBPYxxmqIXyLjRK4aoCBrivK30VCRV8myupPA0Ou95NMUVMBUoikgL+
RcaQlt3Uo6dgbxYHzBFhRwCMwlaxDktdHKTQeulYryyq4clC/rxDzz5ztHnHSLeM
wOYH3bPXtiNdMTBAvU2/VcvyTYgIGbRytErZ8SYk0PcT62mUIrVzFJdO9aZ9aoV9
U14RxMDvdNZ7PSpHuJrBAQ6QUCtQe2EO2jQ/3oapBwIhg14luBYaMpcTCcrBhzhM
flJGIVA/mhn5XBC9TjBarO1J7ho9aas5bIM1aaWR74/fKtYEbiIkxqjiOivaro5c
tOE9shdchpVMt7lzoWI2AgmXkZfGb+B4RIGw6T2AOPGEMcDLVGw6FegkHtZw4vsH
4D4q0ympzTc09UdBlnuW1sQZw80WVzbhLriWGSZQocYUGFhAuX0qs5m8JNJKV2zy
SXU12MsO9jVV/nSKw++WOO2+EZh/GE1irAZZOcgrW2iBOfnHav28oHCr9yTo0649
rwqynfY2dyBDrU8yvPJBFW36COVRTDYbdaNZlNHdVWkqh1YnEP0Kj6WUi9mhjD6w
dew+EuRFOPNFvvRE4DbaIj9o4yRPSc4hMoEQi5jaAO3nw1Uzcv/RFnMxfGDRP4SW
23J1Q99KG1Xxy841yc9dNOSYLFVWqUMWxSi3YUfexcCVE7Ug9pJBflPfUZsh7NFK
b/1aoByJSAEGn2jijDSGHkVJ30793mhEwQFQ6Nv1m7as+cIKUqZfUYTTVIwYb4K6
SyR/GsxDFv9GPpNsYnDVgpb2UT2jaDCgBgnnb5NqBi3/u03uGJog52A+TulgwU3L
jrlVrdRseZCBoHfv2miHScu2UMSkK+K24pH1XDKGMkfUGsyAhqLFGmBWUZ00FNuu
oyC4Isv5Q1gmurJNqe8+jFm/o1CLGfQLAzZ6NxS6ZMl+ac7GFIp7w0p8uXMQ71zm
NSmcaY9889ybd7wwNg/alfMV+qd2r6OJuLyKMoJeWj7PMPPpUVdjzVOBWspvT8ts
HSXBU2duEX1i2B9rPoQvd94pq1FkIwONBfRQVqELbU4GZulT6ksN6PfzZ9uhcyg+
OrEbYO8GPVqHRMhnAJjcRw9aaqRdeZBj3+t42g8cv04EaXb3fwIUzh62b8WsF3dj
0ef0QbXgrE0plD7sRxOizVcrWDy5wwdvMCo6jlVxuhPVGC9GtgA5bo6DUJZt1so5
17vIJ/tl2K4sL4xoO9IWrRKlmrLKdDRs5aaMZNfgD9KcDDBWjyNNoIk60ujs+c1I
vbuc7i+l7uQGwAyd73Ccw9uAVbdYTyFTR+iuInTZmrTSdDrZWMg+v5pHGYu3fJGH
HFe6bi2c/o3+xxr2e1DlQEFggOm5OPyNnDasq/WvGjbLUG38BQEmBXl6+lAmV2hN
sRoG3fVfE0dMF+/MUBqQcgWgcKYyHMhyzC9HBYTp6gKMqInahcyD+yY9IfIOZQN5
Bb1Lif3RyaOW/F43pZ9YSlZH8gsjEXNYEQGtp2KFebeVfLubBT2qv04XaoRHz6RZ
Cwj/UiVLoLSlOZ7UG1pBKBkYP/8PSipIjfYCH19ZUFxyNpT81IqN5c1wBw9irxdu
fQOXhqZMcTXV7tS/Fj5kZBS+kavWq5LHuzUxMlC0UU10V+tkjD2/ob2o6fOgGmhu
Mj8Jn89qhRLrGbc2LyHwn380+jMTGeEIx0T2UP1Kr/Pi6jM2Lf5I85hAA99ZSxSH
jlvGQ0ucvjQDpsJbu3OHTiKR1GDSvp025yF95g1V3MP5Q6Obc6Dnd7upprSmoVMd
dGmthq/cS3UJ8A357VtSLnb7fq2Mx5geUvOlmPM//7jfmEwEYhkaz/dnW+yVUio9
6WiFejBC8PkW0NwRxo6tcXRu9AzHW8nrVNEcngqymOdy4TnQNAcEV45V/FzZ35HK
/YDXxKyV5oVGSHCGHcJbwZ1/UxYRzh5sS9mBgu4z44jNPdigQFQgGR9d3HOorCUp
sohlaYan694ikagrl9HpwmtXp/pUsfgf85j1YAHyXYyLxHT/yGs8LLzKAAQHhNUw
s3/aNoM8SIbpjkfxbA5XXIrpHUv9uuahmcFCaTjrSYR0iMjM+RAne0CKnVs5YKvm
1DZ3d38melnzxExbEtrl2kwYCW2Q2ozb05x/6076fV4etPj8LtXC68fd9sHtgoOt
tyle/Hd/tKJ8w6iYMCpJ/Oe9Mu52LFmLz1aEETAyHoHA1Gixzart/H3C8wy7rnZ/
UGAOS0Zp5p6ksOjLFHVDCz9M46YEXlpQW/nVNWlyiHeRawJ9yv4IBo4C1x+66nFh
gwis2PV5lqlZBA5b2p7YZ7VApCVqvEBAh53ICZHZtLgm2kYD23F6KLpZ0wCfQ+7A
Ki3ccRukE+ADHg0kboQquO1Gapyo2AUgv5ckSrdaBtgLuXGgSGjFtaEJchcRrm1/
oOMLWnfrsLdIy5JZZ5o/5RvAmUBdkjAJ1rh3TFgyIFl/ra6aAENICvRWld0sA261
oWvfYj7eVsMHdm8i/p/8TCoaywJ3L0LbJ2Qb2cmV2Fw/wxEZRu8atOr9gehozLdn
CDAhLqhYad3Ta6r8kxo3sZ9+EeaTUnoIxb7sYXnk8XQ75kz9awP0ygbKf35LEt0t
a9Z5zYnZr8lDGh3ygad4bkOrH6iUhxEdQyQRKDIbRtcDTTgaXkAnRstz9hUowB5d
h/nHQ+Mat+pTu4NfIhkJIMDVPnDcRd2wQ3cmVsH5VVrtkiJb74e8gUMyQYJlZ6T+
yykXYog69JtMGVquhQOxx6t7cJp7Yj5DE/7fCvOxzu2XqT6Bwcuyvdci6pXwXdRM
C7uJBwQSV6zhEvs1qIo/UcfCI8TONkyTPyPArDLQLtvdjDHvhq+T2w0o49cVANsT
T2dnM889dTlBWFNTDpFnnV2FFHBCNAS1+FsOfMMnj06EVChp5u1C+yedK5QiHcsY
Icol7Fq5PfILlBNJvUBfjxMW3YJpBlK0QbFcjSlO+zHALUodM5ISE+3GuMxzxfam
CD9qjhPSCYWSFw88fJKHHKkz9zt7GGahY5M9kuK3E40RInqmNEjMMmMecSJ7aqda
IItaxSqjpsDOPHHxYxvZlqO48/bgTkXUrXfDtk+yYd+StRBdLB1z/ffmSU2WDo1x
ttmiU4jup+vocf/HN4zfZfkLeP9Obwvh5Wl0+g6PyeJI+muPUrOphe/y6lnW9acS
lgy3/PJzs3e7VWh1QSFTExdUvvgYkhAL9mIF9fNQTPxQhq8YmCTSdBYOvJjNU74T
S58F8Ox97eGlQZSSUEHwf+hb8DvlZ5aU5pdXe/IeH9yokk2ymVPzUK8i78+x7/SF
nOe7PyPxq8LVspbsvBJayQ4CFSYiCmqFK+uBybd5MemadsTHAGm+w5t/oF2CDN+Z
vuHZpbpG7rNYRj3uCaSY9ELWfWXuCMjYHowJmh19wo+e+XvBVoogBkW0o2JsHP0M
5aMEHTlYc0j0PuOdKRknwk7ImC/DANCu2UoLgRfCKT9ShV5dNI9pDOQjNIoz6fvu
we/rCYfI91WHA7sCiaUJfBJuKRyotdMqETG0PZ5uGCWDsQ66Crq4WOcj5FYN27xG
sF9j4k0bsNOmh7V81R/zBBeMS0ZL4E4dLf5AbxrQYKTX7ibqN6iphpT0OFHmAtmr
zapNl0rdnNJnAGLAHNa8CyMNdKTv6welAI2aMXBvMGXN9Ex+QpJaWlKE7ToxxNkp
5Rv5XpF6y4OQ8zWW9MTPn/eaJwHv0y1BG9lIW8vLWPgXxbN2P9om3DovB1VVFdg6
J42WV2+jll8uqymisi5XHaHhRH7p1GKmNsp/wSn2v6aGfyKxEB49h2QqLdojpvmq
gPMHIAmptAqrPxRm6XTli85IwNMCGcO7CNpTGl1uIkwuEvZdfpfY8ZWgPNtIrLxH
CzobkJcul3ZwpwD46a+X7Dfr9x/Vhj7ZSCulk3JdMommW7ILJ/Qi2DRyF9Qau9Y0
vjVnEEOQa88BUFeokrfpxay0UMMHzkBHgkCAnG2KBGLrI278qAU8FU6bp3JOzymR
rfZG3CAWwz8fWYNGDFFt9y9X01VNnw3csNQ8h1XqYLYsb0whPgEcbDbP9He8DUOv
zmehVr0PfpY/DUoc9rrX12AxhfM8SALrp4a6s28AxbHdokZtYqgHnmNZRF2ygOE7
0IxWkauUQM3haDoeG+iigbRSV74bn4NN1Vsw9lLJLaDFndqzNtjp04C0TZCOIw26
rkhG5GoW4lYE+oDOn5WNTq/z39MGt4YAw8qOduk1Gltu9JkFQKwNX3ut2qUhH96R
mFPsfWTUfYQlTxb6B8xXDMcQhJ2KdbInsUjFzPZlKVj5RIyo7azfQcSQeR0Z8Itz
zCC2N5Zx5/rgEjpf9Tg5uLuQxBAP84LVdUmKNHBWL3Ms0w8G+xoQyk3Z0otJlBqp
iz3ETHgyJ2M4KUoY1T3w9wB7sUH4NlpqZimvDuL2rnmKOG9G5i1Ka58ljBWckAww
148g+pmh9aIoOw/DuH5KFrR+e/nuhzWOQUX3vY7nMij1CnPGBWz2kkXVUvkEZAic
8z8G3UX2el1FTZLkOWO5xC22lUP5CsiV0r2cJBtw8CSIFhI9X5oStp+eZlk4Tyw7
xW3F6OFbC6XZdWoCxwAYFV8II2TIENjOdvW7mzucRCp2zC2ZZAeu3q9e24BRBKHm
x1a2TVyyjhQZMI+DtF7Rs/DtHXJgZ6JbQDblHDK0L1P8PVt08+whywJcs5Ba/kN7
BbGCSSpHv2O7HTgt2jONQ9MO+mTpoYWtDHUN3HGfBmOYWdrmCEJ8ityIWp1gYkzy
JHJvI8tE6+3qcTR7HJcDgSAfXC7X5IYUplPeVXUDyNYYY5OCbDAnUtoKWxmWqovQ
Pm9BH66WJz/8pdiXolLCb4bsk/pWCY0kGXFCmIaDA6tXzyQry3uk0OIa6VRW0iU2
Q8ZYfnPG2jy8FUXvctiSWrWyucC0/sRa4SdAbhbDV3nUzi3ctHIcTonrgS7kmNIM
mLhx+f0YsXUWHNjAKG5CU337uRiA2jORFlKMAYHNg2yr0ngYgA/WQr0YbulP6JkF
Qd7tfX/krJdGDu7efvrwN66YANa+8hdiFPBTo+jf7jazvatdKlfGzvIh8Ijb5UGl
ovjK7oqcndZJF4OED0FeeJurjKvA/lYYRuAUWGKZwX5yudjQdfImUqtFHDyoISU2
cgDZOyq2LkK0dT51Tyv+bb6410uUGJpbDnbJX5bDNOJuvne1IJ8YoOEe2saCHoJh
0/aL7ph1i50IZcyKH3ED73ZvJ4sMK/t4dAnDn7OahSBrRc/sWcYhyFsQL9bXoe8P
ATVdnSRoK42IdDeJSonWFpuX3t62tAObXyczuSCTs4SI+XYLVGOA40mkDUKhWZUr
4bS42lvYhgBZGBMCqJijv9Aall1tRe0g9GEE7sSDCBOOG0VD9JujjJ3hSBnI5uNF
tEKq8g/VyqBz0bzFCjIn+92xNUc/RDAKLe5ldfFGs2TQauO2OBaFXs5gisorhUMK
wLM84TqwdAlCil0l41v34UhFm/1XXaR+LZtql3kk3jLSLBoOAiBJEaCoVhab0i0X
MiqsvgszLjXCtNLEKe1oSdOtaWp9MXUYIu3nS3pt8j3aOEm+ZuLx6giDuHJb8k3B
eIEA+GfPE219Wc6Jht3H5RZy+w9GBRSfUiZie005DqyclV65UstzaKkbsoFa0SXJ
PnhAP7IiQ/8NI1JuLfLuB0hdpGkU8a3F6GkyjusNdUE55ORPRc/OAtcXlGoUi5nf
9UhKD9koyrU/tAQPt70BpFlFOCMYUkHzI2Q0V3JqA5xS/EIy7wWVJSL2udANj0eY
35hVBnU3mAT0UKjxW5p36/SILxa8UdZmAtMyUG0RBFBUzBetEQNu2PFOKUMwRpKB
Rt7nYmjdNFfT1U4YuWb6pR7MMG/lxkhh/HuEWGVUw03zvrE8TQM2a+A7VU6wW8At
SC57DbQGoBEpPgSwwH4Ladz2o6pFvImfyU/vhgVIxOoJt/rUwbWVVIuA5nX2mGvJ
HWmR3oKshEDzVn42dL97N0taSkNo5ciydikkBUkw/96HtzF6VDzRHLdrFxjfGpNI
aTMt6/i9uSep0Z5PZihIhINpLRk4awvDa5SXaQZR9dz+ubfmNoE/kvJo1YYA1QZN
Zz8MR9ONPuDlRiD8wcqu35G2iheW5m31xdWEbLekMpN96pUiopD5GXw/u3EZeN57
5b+cUYzua8MzizOGpTBprVwwJ9YWuBWjTRnYHSyhYuxcJ67B6BPKyaTbCwly1HSZ
NrhVJIyzEINTVJYm/6yoOaF0xxsy7kTXzJfS1HOwEIIsZOgc0p+bAlStVhBS7k1E
fiucYHTBK7DivICwNLL6kksULauEWzyQdBsfJJn0RYOphpOHvDF/OSTUkTUO0ysj
v/e4lbRda49TRBAbHxGSkgK/pNkfcnWweqqXIJahtXngo13Sgx4dIn4R3RcRxCrQ
V4xtignS6j4r1oqKzz3JNVIzfOoJRYsOeWjkaA2KtyZ79pPchlgfzkev3AAZz4hx
R64Oa+111me9xqNa6gqs/g16DVYqViu9/MY9IX2hu0hYGyXCNh0rb08ToFh3G0h7
yEFwTdfTsV3t43LBsy1QcU8x3CPM6TwNZRo7FVwtBHoj7i0v0+wQG4WkrC9ScjCR
LekY1jOZveUbh+TGxpPn7Rul/fwKJc6L5cCeTsgxQkfWxlqtrD2yKkrtQJxRPm5S
6pGJ88WgumRIoixXERuDqoSJ6KVEgDPZqjPB7mVh1gwt1htrPiilI+8dn4RwlQfe
TeDV4fdp16f+MhvUfTSgLZgnrLK3Lar0VV2weZQlPcacyfmJGfM2zM/GsdYT/fBj
dDFcmccaDv3Ucibpw1StHu1ZgovCx3f6DdNq+gbg2p06xrncKKfg+uY7WZFfDttN
VkZlXMmzJLXtSI65PHK/4fHMN0kuQ4DMjU6H5N3rCtNPeNcGnrxIUFpzJjnY1hBI
f/9QLGmZ920uWsoTWpTSEEMto7gziKT3oGvUmf0T5tMg8QAeFQ5v0xwaGtKYgqfz
3MWJm3o6jTz8vja3tZOuH9G7mZw3A2v16iiKVJBCExpnCwwYWvjKBxsY1bz6NJLu
s0Yzso4TxAqpJ6qZKun5C1PVbKtQjbdoDMWJ5trM2s9o9K/VUNLQFzCCw/TPntlQ
eqNAr2e3WkpvXTOJtk+tFHitXMPgDapR9e9+we+IXC2Z6qpDd7RtaT0oScRbg9qF
ggevDd69thNBagurPgmlbCYTmUGSNeMtW8eXPY8y+azfzGLvjHeVA5Sde9VGM9OT
UcVZi/+HNyIPTYzI0CDExQ6DIB0Y/Ex/DwfH+70cG9a4EIBWXk0rsi+vbOWCIh0i
PhavxqIQh5oOViA1W1YEb7mUwiRNJZqMgSOri21EnMWe0ks7ieNPEzyNaoso9kjK
UgDPwN/rt8Z395CyTUmT25K4Mr4HODsQRQuDi4f9an01aqDPbGuCQxNnGFL1bsN3
WqTqLVNb6I597C95Lo8dufa8Pb97BDpMW355HUDMaEwnwvUZdsYL9il8sn9m2dgi
pl14eKFazAmUgwJkMf1dbP1GFu/cakUH8/YuKH0bTsAujJ2Px3z4xOK4Q9350U0+
VXdAnQ9vA0XH+1sPIcNSfG49BEHi1uqHm8yuyE5AJlfohWc7NBkd1BAMqI4XxR7u
wt05dzkTvfJa/yOdoHxvLwNPd3/m/XPSt8vbqeH2XyLY2LKHS9Flm2kMLuiWZgAe
K7Uou4scjLexvJ4gn5Zo5DF/VKZ/KUAlydX/+HKXJ6tVe47hEoN/1V50PYMT3WYK
E9Savzu4y0NAzFKUPOSVaqjgJr1iaH2A+JxFMChVFHoBK6Z0XbPvv9ogZC979TLK
/Q3SU7C8/d3Pi7Qo7hyh9MjqfYpyq8PkTxdEhU3E7Cals1SCGmvACSkoa1i2mBzr
L+ExPu5bpHR7vCLvcC+TwxM8M+ZJ+euu2wvZZjGYKf1jc2KPkk7KpUGkl6M630bT
ezsrFIdo9idlJv5RbOuSEh8+6cPnEP0kqyDepKquRo8CBiMejSRPn+35x6STmupB
0BqGZxztc+xPTaGkBAhRqsskd1C22KAS3vfG69FaQIhaNBKg7QZ23POY9+VlNkQ6
h8lMvQB6BeruxIs6vSlpJVwCY5znC8F+zMTzYoWhv3SpJ+oxHr+lH4MnzMsVTf1g
lyRCQ5xRp5aK9NiYG7o1UkKh3EYSj/TdF1HarMWAEDKem6yCybJ69DTJc5pfr07e
Ici5w8HK8uH4pHjRKGt998ViivzWjB/1eFs76L/kW/lA5J1hIdcWxxilbsvT+mFE
r/unmA4vX6RsYyjFAp5hia7SmEmSt7UfiSNpz1bEdMcwIzfBmnWBH7vRi21JtjN0
8yxuBmHicqCrbik36N8ulVJZKC9xP6W3skCzH/N+8kPcWQyyfnDz2DK5rxMh0dXF
/Dagj0PU0PKqA9DO6nTCRjTCMhmwzxqGWIcv2fytE+bno0JVFSY6vb67qXz6z3Jc
Fadmsy+1L+5rusn6I97CO7fa3naeENZAKrEv3F6H7znE9BkCUUsLfB+9Z0o91Ax3
QDyaTVnWgFviRLRc3gre4oKfSdVRv70soyqA/hNU3f1RUkVIAzuN5je06VX2jO+H
weOE6TtxJ9l3mpQD93MLUP6ufUoVmaBfU5Py4oztGh0IKlbafSYrMHyz0Olz9JRB
gjJWI2ea4lS2W5sMFA4jEt8ZZxeFN0+05hfAMPqKapNElxrGEP8MpKzkJDWtHwBF
k5tsAjKJsANX4hboBjEPn4YlEEYDYrfW1jnN+1/IMS/aD+SuXcddbjBl9/+HkQon
8Bok1LD2rswVfHYKQH5rmmcyJx4JvXoUTzJHI8Q84ZZd7FYRmISKIyqJJ/q6VelR
NTkl/vnllFoCOs2aIPHlMOFzoeC5a1R0HgJyirQypRfhcAS+Tb1zAB1hTlULXp8e
IN0fD+bPSVHkEXszIPb9DbwNz5Sab0AkFeVTBPdiFbu9a9fLtM2Y2adXu5NgMYt1
Ii0mkksiUXliYAkqtAN25s6MtN1l0+Wl1zCBumazF4OvsOwudPMgNwnu4lahOYaU
GDOyKwMvvjL3i0nQG/uPzPx2pmiAq8BjZaHkotQ0c87w1qktRr2GVvYWgN2vYANO
QRNaIuYQyigh2sIPJeuisfItmKhpbdb903K/04TsLG62Ar/41hz0bSyLOfKdIj4f
LADKo47IgpI7+BjGLqVcabkq85h1XLiiLkyFG4+KkoUOqIij4qmQGviHu6Ji2rvD
3xWiaqf1TIaFJGilZrB/2zjqNfzQ4wi1So/CGffBe4k5SEBJDOInOhk3buUR6i65
MGP9xRuhU6j6f9N3srhT2N1Y3h8xV2X8hfUZHLfpltgffN0JD/T0do3BOn3Bhn4q
OBqFtMLXA0tCHIEOOo/T5aMrXyB4+/gVoCzGgQzspbrOUtg2o1YORpSXY9Z1hioB
Q/Npt4L38L5O69GUcqVJXPosuKmyvWYM0WA5RRaO4pmNWxe5aFCEbjT+X055X4M7
1+hzqRsVdFNk0PcptensvCiiLjbp1KC6qnaDc2VgcX12ER3H5jOGKNjfQloeo7/U
6HzY/ITyyc0zmKkMDyHemp2zrLYsyE8aTCcQGtw5654ps5tH62zhJE6x0X/rGzeS
/0tqKXju1MablB2PhMLkyFcQBVRbRXpo+ePRdcYekKZZ/hist6SoRfDfQNgn5RzK
mCFCG+mDBfpye/Hcv7GdIJ/Uo/zKpabVdninbX2OBu+kgf0TlWWSAe3Pwmrw697k
sJvkD7zkg9uZV5Y+HJCvao7HBCM4bITcoEIxEdnYOmEanihL7ApwYibGwU3q5x8O
C8rfbTHwuUv/Wm1ULx0C3bwwfoSkN9wbYsIAObjx0cJcA7ENmCl6KxFIeHlI8srC
+re+qAgfrVh2LomOL5qeQxvt0mL3Yf6PlYfBODZHvSy/CjX8fT4etIYNH0aAJ0vz
Hs6zHjRDmIAc0qAZAe4dJrocca6YlAvGtlhjHUJe0oIR1HGupAduGBN5nHwHqcSl
f2uVLptdbUD5TyywNz1jCtk+sp6dIf9Z1+qL6M+2cbv8JmrVPohIsjmmkPSMTUn8
J8nofm2A37gmb9tCyb9UUL31AB52j9VHdhoOA/Iio3dAzNJR+sZpLD4nSUyaIUOC
ZriHKSYIKgBQJS7PN4mm8CHsiW8cAR8rOeYAMe17GOBHatSWWt71JbgcG+qzCb1J
Wn578mBVOvm/KbaEiHNwQELsWQvtmMPhdAJBBX0cvkZi3+lJREI3g12XwqVIixaF
K5858u7JgWWLdz37/fsx9jtk9sHwdxVUQWVUYrP5Jzep68dKI3uhyQuJ1G64lfHP
ZWeup0SViPjOepqKPf+baE8hYtiDSNDFHD+URNzs23/+PcweTX8xWATipLPrbK9X
mkHATaUvwtAqu8TqQw4KHl9E985vvBb322BL9ZSCh7H3cbEmmZqOLG2hqkPsUrY2
N3extec/W18+OegQeWN9zSq9r1gKXDm51fAwymrUYsXTdAJ4lgl5KB0L0baCj1hk
n9kXKsIq6yzrnwEJ7CJnZ2drfrPo3WuEUhkLowTjPEAR/NZ51asFIKiB3bs4NnwR
KbzlSLsBjXDdsb+pLGMnDfkw1y7iCmkEN/kSVNziX2y1/VypiiJL6lhJKPRkLP00
AloXfeKvPGrfkTSC811ynIrxryV7n3PTobwR3ItyguYwfPDzA1+Wo7yY674xzhCQ
NzE+AVqB+4ZtvkURto/0h5XxuaSHbmnSVv0sL+M/OmF73gB5vu4xlDFn8X/uF0q4
sgbwUXW8AB5jjzqiIjP/kp/s7NPUJ4DPTQ6j65ffc7AogZe/1wtW3qmhmDaDz1or
rSuaZuPyL3tTg4cL4yU4mEZWDUP3qXdyeNNxG/LngoH9UElq1CBQ/a9VVrn1iGj+
Xj0YYd4PWkb7xOkTtZfIpiQj+dDB8U/bfm/MdwkisXyGzH7vpmJBPUDjUtlyf+b+
g7y2qKwHzn188u1H8KssWBQ6Ll04WS8SqoDnTQMzZrxEwlk9T3ABT7dTDj9Cn0de
0fU/ai/iOw1OFYlmyAoDwtnsaCEsz6yVZzOrWqTG/NFqUPBw6xsQPYTjaxQF1Cp6
i38cAqT0Y1YCyrSKGJi34rNC1yjcsxRTuQVB1ZJWgFAKLn5WdMUC+ntBlZK2csbS
zAuiYi56ChoTqMOLmz5jk4BOVIfn5beOP7RnbC/fvKs29juATPXciancXS90RIVw
DHy/xQsQQTma5cBCGEgLG5q310QbqQKKUlUIICB5Ejh6fclT4syfgyMh2iCWdKxw
coS0itDIdWpWhStc6iGwxNxBmZzFkmWP3zLJ1+nj4k27XrWFMq6Ok6+aVjkSC3hD
YonckfXYtYSEBX63B4pV7HJbXlanF4YZdzyyy/1iGKqj0IR8OP/zYKsRWsL903zz
SZ2pyPuUb44CibzzPLhZ+WuKcYMPgTy2yif9BLdDziLXhrXTgjcplPeoLyOaRt4W
Hn/K2MTu7TD7CWNisQuRkJyrvPrUO7FZgOMjCqiNJYNuSifRvbbPE2QxTcJAJzaT
gUcF/pyDFJalN3uKOgDE4GdheYF0o15lF7CtBC7eSbtYSYscqIYzncw7vlfs+rx9
x9ms03UTfNoAmut9PI72+OWy0KZEohoI1US+NbDhiI1XEMcLynvi1VlBlHBDmSsk
SQDmgTKOjno8gB9JMsS6znI6e3a/64XrGgbeRLhIt7ateWoftXDLi7020IrLTTLW
BZYsCO9cXoPr0QlmF0GNnHbRRRJKO5GLabEffpCRVkpnhyDeCobfXAwtmKvYojEh
B5klYO5GZ/iQpHiUK4g7uX/qIyAF54iARcsYBbOFdUf+syzhdW3ryRJtDLMOedIr
3MPEDWs92EOZJbuYRTeDVowwwpD+W92xEUu0fqwxoPbC1sGkuUcTHE62g9DR+Gz0
8lWcG6LS8EXYI5xqafwcsttSfPsHphXMc1/Wwp7rKxpKWQFODQH8mI9Gd6Vahuag
`pragma protect end_protected
