// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:48 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
RQUkhU+v1qwbf1LqhveXgJZTgC/LJi1RYS4vrjNbwi08qQ4ZjQyeAj61nMa12Lrn
GRFAX4V4UbHiowHQl4UpWBPVoSFX2rScVchQKX1e7YYlQKF/XIhiTW3p5GM9c4en
SroxILA1eRbAI5q+DxaNuOKNRnu4eE/2ffGtxWXFSIc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 2448)
uoVqU8ZxzS9EQk5wbNer2fy8cTD7faJCd88NMXuD72ND9WBiQTfeumouQyiiWddF
pQfenIpcLUilbFmR/0BiS1huigMm9eQJaSrPOZiMYps4VyBFeFy9ZdmvRRUHyocl
ZhrGHNJoWTToE8w5bC+dp5c65rwJCva7YZGYDrGeQDB2BQXR446sEXFDJU1aEzHk
IjNiF54IEBSfUqc4Wh9/ia6tfiFGEbIyia4ZcIX1gYo+8kyb3zah5AS1UHpBG6GQ
FK3ViMEGpcLGkVJIYO6t5qMNiAg5nGQ5C3d7xws5v5jmd2jnbvXydq/1BucAakH/
l3wmzMF0Y42mKHgRehONF2YJTga9rb1DFq/AkQ7wHaQL9PcWWLMnbj/X2TOlxHAm
jWIGx6EV+wUExZnDted1F1Ejqt2ljA+OFIXkFdFqB5+4RECPSP1RxjFTNP4cR0fc
vCqTDpOfFPfPjDM00x7IhZOWsifj0pVZxv+WICZqNabX7zZwik+fLHGZdxjSMHCI
unsQ3vK0TKuclYXVefY+XBJsaw3fwU4kSCXoxMXe4uaBIyK0UEoizt0ZrqpMS4Bj
gobeIEMG/vyE0I8+SadQOu75O8BnplZn2ZPqwewdKXxAOPI5MhiTZTCq65c7Ci4m
2AgwRCvcMEKmb2klB6p5HCk5UZOcWhOqsjIrNHvqkBNc96OxNq4RNYavRD24Zxbq
ASbjYVmAm+WbjKB0qOXZ9r9nM+mSQDtYoFf8XAonYgjq8V6+xBuq+xZiG1Bxwpu7
Efs28/5Ahydmq4CPDB73xI+WdKJUVGDIsXMWlWdgwRrO6ilbxlyn5KZv4MhgJVCc
V48KI4JIKtw389ve/0BIKR+GMxm7RbIAH7eqwgs7PWfpo7a3boNxIF+M9RVxvgJC
tUfMVlkFQFx8DoEt3rMN8dKFlnmcgLhzTWEeI55nxYZsb7MlN8SvQFF+13aS7sac
EWu9CykuqA72htJJFOxTR+39J5zT544qnAPALyKXOOzL0JadauQlkJvMIzGD5Mb7
6+Wx7RGF/rQtAbwxBbd7vuNJMrW4jczusVkKUDFZqLT2H0Hfg/oPwzuxhoA2yjft
6okxeiZ2Zp5HR1B5wV5sG2NnHYZJ3uxu7AXYrC6DoxEq8Eyb4LAk7LBNkxvLoEfA
UfrUxrDRCr1xbxIBVou70t1GSfJnnee5v96L9i0W3BID5wha36wolyc8FNDvp5/4
pKSvAvRjJwE8R3L2DKqij9kZAY4sgGI3JSDzcen31EfeBka9U3yLVm2g+lZAp0cd
6f1YdNgaqcJnEDRgaAwgvgagXSRRFPaC1ZFWT34o/BEGHdFh9SC0ubZgX+8KJF04
xf2k/jfdtBnr9QPxozSxp4JPDwXgdnhUKWKAKeWufy50mwrOexzpC/XZQPgQ9VFt
UwY2sPs69SA1WE+EUvUvlMa/rc7d2fT4cjRdm23Vb5LQX93mMJn9PdZl8WxY6ZWF
pkBV1EpU7cRXNcDhI2FvgG4N8egvwkScKo806rf6k7+Zx2GmOmYsIBdtW+/H93xj
ljdh/OCq979YLt+cYh5QuUVoSkLTX7zmVhRInFbjHdHquworAsfXYFv+I+LWEH3t
Vht52sgdyZJ84hsmDNXx7qyDKGzSIiahhTzxVx749NeAeZ21mat5NjVh313pcV8N
nyvci4LC/G+Ok9jqDnpNZaJjDo9J67jiI1Wd8vGl6hEa7obtJeTZtVEAhC0yadms
nnzbg9py5M3I7aK7X/jK8HMa1o58wau4BXjWE1QOTv+Ar6PY3i1K/nzxAgNi94if
MCokJ51t7yUPZEx2YqDQP/6RGwLEAssQbMvrLYCHURsygOORzyMA011+QX7ogz4+
UpiBTItqAWQTytJ4rQA6pK71NbL9Gpyx7Z76ALfQ59ullMjVt7bfq8qWITsXpVrq
mlDlG3YRrT66E9MNpatJPKDQm/rCf4tBSWJjyLtpv1dkdK2kr8fRSqW1bAnMcM3b
3bZt4el2Tf/+AIL+DhQ5Y26mk145nXRZtKMYiHs22HqfLA4RE5NjcwdpKJPRbDfL
4ypkC2GIyV8YXC+hx02Pd3Aexw1AXU0rtUyATa+tjoVXo94M2HHUAnjh2Cw2Cg/p
XpcH7KJwoHC6dYdQabiyF7c0Raw6bhSFygZER4rsfeIkrhQe1JhP7GQhGscNKc8O
M03u4Tyyk6T1qP1WYnY9LwaPQtKalmT2DJPbA6v1n4ZIoW9bOD12KsfawqSAIQfy
iXMkJLuy4FoVdPmKIXQMECwSZ4YeWn1BCw5wRxhGFiyuB9r5bf0Q0xYnwbrXnZnP
dZ6KlDTDg2xOxe9hJHfH3PEk2UwRSsqCupEOosqKxtvaBrJ6u/Mvl4XjgAdmTgba
gDdtRKoUrTApmFvPvgSpbS7zybIun1Trnh21v6Ugj5Az+PK6m36o7HsPrhbnRu0A
MfowNqUEUK2xcBZO9YCs83su3snjdQSuu1tInzVmR3sMrU2CYn2jWsV5NGyOrnbV
Mpv+KBVPNctob93vaa4J92Yo6PrZQzDuzk1I48+wVQodNuTKBo/XUsdmg7IZ8nhu
igR1w1+m2CqY76KrYd6HeQAxKB3FNItr5LzVyVJ4UGFIY84pPHMqGsgDHDij78QW
RL6fp8hxRgRjPzjJZ7RKJWhAK1sW6oGr7HaIY95fYo4zEC5EtzEBXoPGDL9woY7x
wU/4UzSTGh3+yOnHsqdaNr7W5XrHVMHXEFglGf8UO7U3W/5ON9s7YwuNA2qSxyoQ
FfsaqNBANa+Mai5xKoTcF3+SeXV/D3ayqXBAQICBfQCDqO/A3fPDnw+62+B6wbEW
h/gBCsySTHsDgforqPsIHlSg98iPVtlRESnOVE0LJFlbiXnuJ9d75musjAnYirUI
c9zqimI1bi1YROKfyAVLjU+yKFYawhfr+7HXjVQgZvOp93NNoBelC79PSYfkwzrG
AhWotKuvg7rvQt7PSdcD9aZk2FVUZ+opxdTZyYrKVyRahfkN+kPtrgvhPSfAQazl
NigDn1hEvX66tp9yhCblMFG28XfxAnNu+CAClf2PzQGAyCJ7+FUglZ/v8RFBnIX6
rjgpldpf7WnaJZyLsmA5DyUwt0lxt6oRfVvhdiUwZvm9m/sF/x67NIfcbPpx0WHD
BzrneXiOB0id/vFuh120E7EyxLnX1AHrKIa7pHZ1kDm4+pDsjmwKA/qYrJfkV8sR
t+/3WuY12bm0hvoQq+17pcZ45jni5T5tijLOIzxgvYeSIkpQXzV7uyor/VKuRXN+
`pragma protect end_protected
