// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:55 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
bCFWpPH8OAnLPjJZq6f6F+hF+bNq0SWG+tA8+L5jBKFhpE6phjv/zxDabuOdBRwG
LamAxrR8yc5JWnqlr9z9cx7mwghV7+hVs4BvfhwNjcfyY+OrT0OjJ0YU0p6cvLXD
lYaBohp/nd5kqOUM+6ji6f5Ix96GWA9u7evT/5o36A4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7328)
p6bqcTUcmAroipI7e1uQqCTh3aPZEQtFBkxB62lMRRPy5YYIvz/xfkahg1z6YiGQ
pAvYSPGMEuU05GgnIw6wg5hg5o7V8mXaX5cy3UzuW3AzyGxO0eudE9cWt0xqOFzD
Xz9bBhBT2j2sMbD6j/C9xF7YJHRd8BGnvlODwfdCsGMSmx223d2eofCbgxq2jw+k
5eMQ2bTA5sIhLL886aGhz+hAv6SRazDrQVPCFEEDmoBhFsshTOSd1tU15vwbwpv3
QHGpQPwvxBH9U0XZAJSDoGaTcYlRvvmsfZEf9hTX9woJdrt5fp26LjythByCBnA3
zQWHVpvSBrDITRpDawaf3o3N1MaNiec6930GQDw/Ko+EjZToKVz8xYEzQWTJNUhc
KY8nsGvl2AZ4T6meIqjxKXR3Bd1WPp2eSZ8t197vvzzHCrsQWl/jx0rNCoZGeqAX
gxz5KdWrtq0e51YHbylM/dnPv6lfotuv6kRwYymKYaQ1EpAbFp/t3++BhP2XlCa3
rLN83hJB0vwHRFmr4WYbKlZIhukK6bN6a4ssl9BsyU2Fc+uS7JAigisyq5unpYn/
Oa05L2SVOZHXkja6JLDajj0kT+WMYYuKVKk6jKsSjPX1ePwabn49rfhxIX2IJzT8
OD6IEtNpekqWHsPbm4gzvwEP0PArhndY6ZpSmNaCInsAg9WZafsuTplOjaOoHzLk
96nAymjqp8l2j7wL5BJc9IFl5BxYWtxc+55np/CUCLa57Zfo+oGu74ys0s2BdEWE
7UjVWMo6m/5OSK6DrmT+S0IdkmN/98BAu6eXXypaqrSBQGp2fRt6GzDTpT519dcC
MPBlOQjUnl2BcOXMQKyLsfbO3vI0gziM0wYFB5F6TkwCkb0g4S3ZHfjyF3Sn+KRp
9i+xTvJQN5hWUyRObPccZBGmOFwXUG8DkdR3njOz69dqyEYRgjm6a5EOLn+gECLU
9aQNNOwaygTmeliou3lt2xLXkjYqPWwpF8V+4e4BZ7xjN/+UB9jd5kuc2m3Otgm3
/DFZFoHAZgLehAkn+ikYWlNdmK3oEK8dk/H25OxnZHO7T7sjvzS9B3U5Es7fZNkx
P8ZQhIPeP+VjIahsZkUlnDiDCeiYHk8qpGrN1hkyb05SZVhvtbzvghz2d9HMNoP0
VrfgJ2JddmrK3YwQjLVgqo9LdFCAD+LSczIGnBwpN01O8DLhnv9NxoNstb+ev9C0
wc7Tc+PNedn18AQ0Dr2XyEeRh6ZtdslsMc+xXCmsqvRR4LZJEigBmIDpzWuUJM8V
dpjxDKxJvT7mPTgUcD94/fIKzez+CQ3LkS4RT4odftZfELvUmnin2qLlh+sAOXa+
5FTSpNPapViwyqbqEmSRIyvsOMB9ZEPMkTOYF/CCF5YpWDWSaGOG/NdKh4NmXEnw
PAUSFzaw+ZVPPZaVgDS2V35RpAIO1JQBSqfelOkAyIrdWAraLylNByPu2guI2ZOV
GB/deQ54857mPhvZ+H0U3bXyQttN6o8G/e2rC/9vvXzvCh9E95bxMS/m7vumUxGU
tNjVSwZHDJp7FN8v5Rd1tHXLWE544N9sTbwYDhYex0oWNxZM7D7tt03Ies8WGi9S
92lvubwfQjWv1gC6dv0Ico8WG1FaI6DwHLyZpuZZ0UoldIPvqwL+5ZmRcL+qD3xx
iijM+15K1JZomvEHKy8NbTyzyfI7/62D66qorZFIxPTtTjbwT/Hv/cn2+ogSom90
cyYJEbG32uybwBSf71iu0hqK7fjSep8ubOY7I1j3jK53xPsp7RxiTv99CDPbDFFv
9FDqy2NQ+feRTWbsBTek9R4evmROs3K28V9qhRYgmruavni48f4jL93Y7H6Q9Ktg
LgH2f4kMg2fT4YQ7GYZvQJNbiOqwvdpR6Zkjhe2QgCKOh7XXuF5nz8By91aPnixB
M13BTncv/8ALk8r3H/b7K4/bEtqnGWje4GxNT3bMBXH0+EmBluK/5gjdRNjgMNOR
z5p0rvOmJqE0vN49SCB6PsrgSVWSjc3E7+cwMfrMUxcUXrLS0aCga3FVtVqKCI0h
iYnmurLJVG1zfXaM+3Cb9wzpmBqRn+GsQkslj878UCHr8qxYhD8KtUT3XfqGoxPB
GGU4IRPyNKjjoftPRH5HuYfTUovI42FjlDMBF2FUVx93/b0ePXcd5u67rhcQSnEC
8iN9ZhqNvYFXQ1BeJgB3zRxR9WII4PuLCRZ7mU0P42HihbN8XV+LGO2cxxuK19rU
6Y1H4y6o4xMkNsyrTs3a3SUDY5//YWSk4C5gqo0y7r8d3YDpY/IqrKGH8UztDeCX
V8mfMLnRmmOFbmdNvzFWUf7IHirwe83DNHBKHQ8ONEiVUmp0j8VsgIH8uecK80Km
8jbVM14oStFtJ+l1JKgYZdeEE+PmbbEUAWKNBAMiZG26GvmXA1blDtJ+iVnF/b8h
/nrAiRQjzQvu7iK/CPBGtbdLvaQhPQlLG2dMKo78SKLjqw6ld4TcshebF9anXUCc
TD39rbm96VHLE03kEboKYsyV0J74sO/q6W7eWT7k6tMRr2Ca/ipEvesqVmW9As0b
Jku9CBbnhixWGOHzBMEHoYzvsUdJykbPIZcBrXeHTJifWjmwSZtBXc0yWQEH/EUE
eNNXB+/y/mwm79mwZxnZSKFG9oBtIhMNQiCxufv6FYSqPqek5M4qxh5o9yz+rBL3
RayEDI/dqVrGO4IJRK1+R6c+33pwDiE8D6iVqq5fyzuRg+Ik/xBfIlRH3Cngh4rm
mY5Q2cHMP93Km94xQbJtzZhkKPNXJOFLodfSmUeaMsDr1oIdmGko+xII26KrhWBX
eviml45W4ugwg0qOgcpltQvBD+GKNSGwxXeinNrK31QZQHRnHrKEackdUGr/qVt4
avVoT8l/SB6nMTwdTixEE4BPKKkYdx+/IzlERrG2uBoNTaQcRUaM9AVL/Wlkrhj4
cWS04ueXcvNS7h/RKoQ68FOqLi3TA9oS7qV1vd+yFk0/1Y4v2gdJJuHs5CBPK7no
+85z74L7WSccgwzR8pufF0LY3bfOtJP/T1lcjnlODOE8ppEhnekN4ZtIrBuRLTuX
DoLYwYKZgVvTWXHGTBEkkLXydudFWALmpn/6UjALsZGQbJykJPAO4ldhdwvzIWMm
kPGjy76DxDu9VRSn1QV7F/7ZJQt3h+/4E+EB9bTD23HcFK6kUalEF27XnCundqWj
6lw0lLk2MyRm2scC61fsvP0UWYw+xGIKYnfvGF7Wqp5DLbW8c3RwkuCnJR56ne0o
4R1PjHLudep7K2mMnPwflc24/T0Aam6iLDQQEUCzYe4kV7pVzB5EoMO6RzmAJcap
9QXq4UoDK7zByr1JQTIYpsBhwLzzYX6eHrCMaHF7Ru+tLdF9cZcRLBpsX6kdZFJO
qy3OgliRn/UpUQO+wIUJtMcYD84bZAjjT1V2INaTmaiFIDvDnuo4jl/DcuXg0HI2
GInJgdt8Uz0HqaI6YCODT3h/0AEUvQlxxTJqKu7+XGRWayFcpbGhNCh/UaSw8Jau
9O3K1vj9LtMiGIaXxbwJSWB0K/mpaX8qo5ngsTs7BYg15CXZ6Dcevv3jp84YKwFq
jiSn/nwJeJPODYaPZzsY3ARyBFcsPPLkUE54/PdvISD/qUVGikIjNCP8HHB8+sp+
OdngvlgXbp2PTK6oZHMYKb2MhmL591lhN/FgyJ8BsO+RrhqOlJtyu3u6AMFk1HlH
bn1ctBZgXD3ayrzmBdBpHjWlIYe31vCiQHhawQxKaAahNpwmqgNK7fgY2dWlphxJ
LzYI3PvEhLyj4zqE/d112ZOkEihx35LA99IiMT6UF102lWUcyre8KGGdQ5vHAZgr
sxq2x0uOV6dgKI7f0A92I4k6yB4qThIMbBhO6cp1OGznM3NEw1A8zuQvEMiAKKyv
Ywuwq8ohfsiykQhq4/fp1ZtrZQ0ZtVckVeMLgP2ltkRKIFkdh1iK1A9eIfHlJbLB
habZssMhRiXR3VPvFNdstYL+5rPHg0UrgEqvBhra/MtOVwzlBL3Hdfs+Zi0AqMnx
/N00g/4FDboK1mY1kj8Cpj1ds7FoXjK9CqNExR6ybKFWhFfB8iygqgoQlu1X7YDK
ltBOlVzEC9euE7JyIr3oPEujC19s3o/YEkIcYqosNZTbsJFhhMmaezp83XzxZw/4
Q9D3lQJdszelIFnFrjKRg6L7Zq9M5mg0PplQE1Uhifx2MVrJkqJBNA6rWo05e/6e
2vNqU/jBYsi5mWlh+zGxySDxdOhE9NXbEPuF1ksmlfFzcuwA3ObEdqKk1HvrrdXs
whdutPrZpqmopmZaA6ndCVDwkOSwQGe6huR/26YYHuhHdWkUAutSr+619IQgJ9rr
En/JVCWFth+CT+YM7afFpdcL77hNIo63HCeluhbv0pFrYUIn7Rz+7pk9XIo1TSVQ
O9tr+ifrRZZivH/tsWArosCpIjOxFIHRzX4+orS9Amre1EF/pcZnekAHfqfAsETK
0z+dYH5M6wJiqR4e+SPh+hdrhPVS1Ea/O+22b9fr91i7a1sRkVEG5FSFKEzKDmuU
rsdFXbi8D1sFykZ+dbixcs8YH142EpYpN/t/FSz4dXDQ60r9g0hf35knk5vJLz2C
DwG/Ez6YwjpYSdbhJ5xAhVJndQUlQFFLEVJufIzcBHSUNntN08j9QB7gp24imq8L
aoSJBVqtg0u6NWV3MNH3rWlMjARNp7F7CSGthmiqCP+D0+DTfQWBcNueFMK/t3rT
zhnTRbxEsRwroUjnxz5wcAZBghJtCUKxjKHe03IAszRuYbT24rYu51IvoI5eM8GX
wPqgFpV0giJfX9PqhS23AD9kbRfA9OSc1OsVCrzgvzAVNYI2kcycNnALPA9KblnX
m0tpR2LGPBDh/0TGdvNMbRZqegMQGBF4j7AOzL0Hg4ETt5+ITp8jvnx5KPu7c/hV
E4/TKZt3qFim68i2aYiwI/IAbuF79gNvmUM8hNCWXwLAz98Or/WmN92n92wLkXO0
TPgoXp6sOZ2aaFH/5fyt5+RdsU8otUMXO5ZNAT3G95ZmvwEoPyJr9/sTiaaxjeMf
ZyfRyD2KOIiygxPzR7Obk24n6p/cMwyzUs3Sv/ZVzhSeOPeUF1pd/taUK2APM0pX
P4PyEFVfrZwV7TnnkJ0FBEAMrIbVsMnotseq1IM69Evoe7j9HbHNBIhhP1LaiAHZ
JlLfVJxGwyhDPAc7E63gUhvp1ggIieiWul9Y7OpobwA5KviafWfgGm1U6CRYolUA
Av9xBLAtjfVPtCFSZnTfSHXxQ+FGlX1ghTAXcQkDbuwkF52j8xOA7/QuxtahB1OA
F3U36jLPYWMtSOwD+wx9EisUEmqyNKoje4uhPxwwJLvWlCTFTuUyDheDTk/2Gfvz
CAgY1WzBe6KFdXuFpTbXpr7JiTnV2LCKHIZ7BPm9RlOuTBbkVTZvYRPhgy1EMjro
cCdkRA9VrBPx4bl80X14nesFXhAVa1Q4e5KYebbGmfm1LG4LOdjHMQheg5jE2Qje
HFl0vKws7sGARUuFYgmSi9hPBQ8KvtQhfyb6TXNv013CM9pgtM3FSRaFnPo6HyVf
Pmk20bubFu9vQW3kptK+4nreaSVF031me4bFzMqRTfrkXjX2cJtq1p9hy94va0Nf
1ACNFAWcHFBAWZsz4uMTEdNeWzv7p2DkpoumUfs0pqmaXUmV5EzLg5U5FaIgH39V
dRKwBDLbt7Z6wCSrJRROu3M3PVTIpTy5gpqfEhK53KCSYb27pwONye1u1bPY8+5p
exCZwhHZaVcUm7tDdR/PQXNOcRLZ7Knx1G1GYrVSnzTq2TXXrHjgn0kSSt2ItIi/
JwaAnv9OtHmXHBAi86enQivb+PvyL1tXe/3qz2cf6gOVaM7Fo5P56Y9Yes4qcC/C
DUh9apZI79juzZCdUz9ARo8dMvrG2NjfKxmO248OGp3Y/pNDlCLmuP85O+V0HfpW
HfSo4zpePeeGRDV7QiUjp1WZGCf0uey9lu7JxQt3oZK1t6NF50HnP1Dr7xjAW+8H
ROs1C3sBqxjH1l312ilOj7yzv71cHIz4fY59LMG2aykTX6aKu9maPDc1IlWLo2a0
14wd7uBS0yTFGXJ6bVh6/3gtBd2XQ/wOAUT0GFAk8zy/xs5LP7LX/1rJyPXi9Th7
SUxl2mYrIW/APqDv0yMtElBvUzaIHakJdd9eCeubYcTWMfgEhpyeCy4cRS771Ajx
ilNFCw8FROV+rMUeS44+aMYzFIa+kkvUSovNuSEQv4JnHfYlDkTNic6CFn7oVK1W
V1sP8OApVjhxqiTqdgRtBhMqjwgn6+dwoyaxXfK+sQ8p4Eji1gkLCisEh0q2JmA0
The/XzaRaoq4XCyDRAhLb+EqCWf7E9oSinPjDGRwEPM5yJ1nlnZU5/xvXg3q+hFv
99laasHeAI62uw8FO4CAUJamDkCTHK4JlN0q+XP7HVbuwsonojK2IWRdAAYv5OcH
s9RiEyiJSwGkGpQYbKMgsNdLIpuOwhRZbQP5e7gtQ+Vg4LkFWtMu0WVXh4/aPIJ+
5578fH5pdpdW+rQOqEMXYV9HBKC8qXrfas8h2bRQgdr9Rmx0KJ47rdLoaIJ+PxgQ
MfztuNguM0M38toJhDZ8vMSsLAfKeoLKg/1ZhN6H+Pa7SEnZkoYNoHu0dCNxUBVu
ofZDsL8MlqIucLHX+vwdIVGRK5700AF4ExwsyJO+f5VMfaj3DSxiIaBvK5bHR/lT
pmTY+TSKEAsJVLfjKLtG9tZaQB6KeU45Rx4gBXNeQEwc/aJrGO9JqZ87g8Xnlpg+
Xv4cHmY1GkjZP6InmhYVzhZ3MBDriB/ev5MciLkoHW+n5UC0JX4tX1gYr8WvC1eZ
PisMEhNx6JvpMAV/npKVnq9ZliIwFTCkuqOFbXSvFM5S4g47vIqLsAP2xjMahLwT
gEyC45m0puEi89BdbOUYf54Axpe8pjSv2gE6+b+/GTLMjWaH0tk+BDMwC+sSrL+P
dTDz8ihvv5+a4muiyKeujhKlOu4Zz+dWgXYbA8clBe1z5WGunuBPd6996tOVS744
qP7zZ4XxgA6+44kMlGxwdOl/DAlRLESm0YMqzhWYj5b/F5bRbe/lHAKQgBDBmVKl
IkuUXWIqjKVZ0t9EleFlhPpJV8V7Ggy33KGGvUc6BNgPHW7FUnRF2QUzp/7piSfS
7dYL3SBw3gcn0uvw7j+Ojt2aw9x4GTeuD+puhqs087sPFb/gTrBAjMtcudB+sVUW
eRfrHYGisds26CQO3yMwfWLhUmTsTqUoXLe+DB7AUK1wVL/8Dqk6pdAVWI14SE17
rv0dhsvYD3vGNoEW5zBFGtozCS/yyTKy5WaRoeSd0prV7Ob55Hylzu5884qyUxef
OEZKKiYwrU9Ol1USlKoKQN00K1TiympMx9oga8JVFb5E59wHDj9np/R03W7LKMUB
br+QHqkEqnsuPTjBqlBIggjRINcgNAziZwZlA6wFRNN0nSyyXXy9qKd/1NQfMI6A
LfAZxdoq5s5us1mP8eu8WvJcBhSh9vPdXjxJ6L9BiSbVfyqbz+RapzQGMffXqiHV
eNzA6iU/lmZXqc/DTcyrxX9gl+KWTpk/0h6oMP08+hRR8j5sS3gzisc7uyN7LwXd
NisQ593DI4RuBHWb5Tp2lcUY8UXnJG73hiH/J6dtDviLrNIDnzScSsxsOwgd+FRi
zKtdTvHY2ZNkbwCHlfkT7lpuDqHuUO2Z8LhKCC0N3PGcVPv2W2DLZAk0ebPBD3le
SMXR4VAeJZ2RkvspYzrqyQOpzpX+Q82dPA01vyo//yaLtExVuY6QP5qIHBALdKv+
ioIEwWSBWLDz/G48PtF53wckFFErwrf4A5oR4WgEI6Ov/GFHOARGQ9hTm1VqaGU6
W/TZXqIoNh0lqZtICOy8gfmRSpUt1X/jzVRL5HLiFVr24KprLMvHv4ujT5xWmq2l
fwtARBRbpoMxSJPyASmZ/cMDBe2EgUtbmVFAamw4BRg7uD+zhieKM2OlZ5GfWPX6
5Odw+lvsPs9oP3gFxTtOjfue0djmVhOsIaVcebONW7e4DP8n26oToNwx918bPD0+
pdOyKWtLBZBtXdwT+EuOJMI2BWw82hkyUeb/Gb0ztatpQPdGCJbTn59BP2bZhqDm
pE/SqDN48gpV0NGjsTf6MAkA/q/erAR/nBU2FbFu4f3Db8hOITBVfvEw84lftOOC
gV06iar60SQ+u3BZYABqdPcN+7iUcU1c1Us2gxl6SKuP4KUNVxkblv6ah+2W95+r
XBioupk1GKeoiZTeNZYXDcWS6D5eaTFSDX2qoNiLZdHPFnoWo2yqL7jAulfDyDZ3
2sTroP2csN6LUJ1137wvhFOlKGes8POvJ+YHo/QUPPdYMsCKVNO5764p8Fcgdq9g
BxtLVGEuugtn/Vm/ayxCHi3+hqv16IxJt2WjqsX6HGkpbkFwVKpMjL2DKHLYl+Ct
o5yMjYvLYbx3yh84RMuHIX/EwgDn0VDe0h4lfRvDAAL59n2Zieh+D4KsZq1oxkya
IUDosWMKCefh3W2qIkZsCeFKDJnsqMM8hWx23AT7q5XLF9n75CqxPzJzxWiVWLcs
ROJ8t6fEzvGXO4g8ts+k32j9xJfmWRGy3sRVizyuIFFOMfSxOTSpIxX92Fxy12cu
D4WotgkbzTdZqCg/TQfE5KnRbU1+bYgXDW14n+ssgaaxQctQrcZXCxH3BlB4nEVh
vLYCspzIMp3InXXIUvJALoZwt+p56n0Az4vxTfSL2zULt2pzTujNJAioAU2R4BbE
0aBXnBJm6Lm6SPS81qi2a5kgnq68N00nJ03sPk3XB82sjOiFd7l/IPa1OnFTR3XJ
JPMVHvnzqf+BOSfCd4yIQeFH6wEvZOapvW5x0C25QZ2+GAaE4CSjwpsbR6rnJjtn
BovGUPoNH+GY4/lcW3gXESDjbg9i36oH8/JmKQzwiCBai3zfCuxz+7zBd09zP/hj
C0iOUqxHKNyk6rTWv3mRf2/JM7lB3HJ4S7AXFcMQzoJl809CpEu7RNVUykixFadO
DpJDHoXcgXuW+atDtkFqw5HAIaDRiPEYZFR61kSuorfpAP84tjnyaExHHGek+zun
0wOKwpcJsPMRQuup/tCFBr4PFb3uwrkZiRKD16LAo03Uup8Y7gJW7VmgvjqW4mSe
TQozQg7zMxacAMDXgHlFWrEMto07dYNXmcnMvREsE2dCOB88CxnFhp15VRpk4YAo
HZovnyZ39gjvuafQ2ngLwEjWx4BQEfz4LG1Cdi2Jn43Ib6GZg/2uNPmerzgFvgax
OeivmvblonewhBgQqwsfZevT0JzzN955GDU2pG6o7BEIesDds2aBx0ztwGUZMohl
zvpVLWgCosfTO2gLcrLeA3LuAZK57O6t6ZgIKskacu87YT3HEhfpgu3SILShICRF
C2L8UyJKoQerENHXCMU04yLhoeAE/5di9tXsIONTzlBIw2VNoNwkY1nZd0wiYKDS
XmnOYxq9tQCDmTFtaCfIB9ihNe/pnHs13aLJsb/FqdopzM1Aqx88WvTgJ/4T8LBe
lXybTs/OWSnDBfN+C1KlX0NBw+GzMr5VwDFCjDMwzXC5vXtMQ0mJwboQipdfylo3
hYnZS+j8JvO7C0h0piaJji7S45dcI4oJc4Ut60H1zPsU7xrmoER8Va5uIGh89zEM
HcVMQElLgoNuz5FmXm7UJ9uzV+gWwWLz4zaLVbdMQGQFqEYXUrpN6sHOsOIIzrli
HZ34pPYdvkMWYtYLh2S96J1Mr60LmoGOQ+A5zLiokC4=
`pragma protect end_protected
