// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:49 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
IAr161qy+G5XCWSgcXlwSvq0DJyfljPTGKEtXF9YWR7sxdTEkJtQRJIJeAfiS5lJ
M3JquZnc7WD7KCvXclWhp5xvjyihooXtrbalsBiz4Oqj14uBLzExqco1jZq4VxH+
sUtsGBgDLvfnFG/uxPVMVS3xZQa3wrkeofGx7ZgC8Ho=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7344)
NA4rc0abcZ79EA+jsXuuIhvBiarQvLXF0hGN0V9skTXf3Oy/SMhHriIb55HzIUA6
p51sQ6oOJvEY3EKXg4SIfwzvV4n/nNGUNcWHStIEral0xqmI6NiSZBUU1H97KYfv
56+pytaBS+mn+6KxtuGYeUSus7caasALfkW5nOrLv7nEpgHjF3F5dHDEa9JK3KJf
Bt4m8CUqB86TYYzaczjnBiODJIRZejuaOqcQE0M2EMWObNsCQXXOFXv9rb5agaIj
MojlLcstZv9dql7cfpiVBvvZfXDZoNPHkgvdo+gqm5lHyaksupGXev+b0QkP6WOU
BeIDKHRuBJzpdD37MEsJcLajehHv5YTUe7qFeWShyoGRLq6/o4q4Iu64G/EvlEpM
2qm63fB0SdKRblreMsTvDUJdIwR7gTJU4DDO3gf/7Kv0rVNBW7asTXnS60ESxJuu
nuyjO8OXa3V8+rhJ4SuoQSKJ8MRzmyOQ3q69g/50wefI4/nRToFid9sQGKKZr0Am
J4h3MsvZ+b6eyunPFp81b1CxeYl2l2qMvHvS7roa0mmkpnI83SbIApWm789izJj1
upKcPfvrhS2toRm+IOBP3MYdWMr1WN0r0ZwJXpE/BWvM7OF6dchaMS5c62/LtZ36
j/T06jLsNqUCp3cgbgGa71KRl6WbXw9jDRQRyEVTvzvPBORUTzGC5VJxyJhvg3Rd
IvH5frfLVvr4YS3rl4SGIMHnltY7ueY0GUvyKAjjlu4M4zu3+IQvrNCpHojCm0LR
cYjLJY/u6RVpwiiIeoLT9PTpvdL7sftF5rl7DiJZYh0KjjmwkANQNSiUexUGzos2
gRSsydxqsQd5zuM+EvnvD9SW7qQzz/EkwPWlDRv70wVa29DaYdpy/1BFjDakWAOD
0LPpB5uKFya3PHfMuIX0zzn9GO/2CUl7COHz2d9GyVs44kKWDXgZ8yxhayxMFIst
+7VHMIqcQGjAuQzPmAUe3GUD33k+ovs8BD72Ewgt+W5YcXOfVL7zW93vOfH7E9bq
HeVTRtIuTotI9fQ3wixB21radwEMKGj9xwIdmxDjD6VEoFoPRbqLIB4X1t0jg8kn
T5rasBJjN5zVNbzvijYZJydZQKwAVgFi7bR+Yje62H1jIdAYL1FUK5GvePQolJC1
HDAcygAGo4L2jikxl72br7J0bH62nSHzeVm3sIMZsaFj46fjIGDocoI3IJ5iP1q7
fO6QBNqd40OWAqOJwCksFxyQ+Iq2bzdSFbfQAuP/9Q9M1q/2wF6L1U9EKnM5cx7B
+o7V4Rrh5kp8lbd0Rtp9lvThNVXX+4l6jL8OTomxws6TyjkfHbmY/d0PH+/czKOb
yGElrxrj1AokdU97baimzdDgz2E3MlvoUMHHd9gwUEH6KCa6EuFFMvNVKxXXI/Mv
5Tzc4RbQ0J0GK7CUbOUUmVQWInZz+W2iscbBNnTvk3b32QyYB/vpL4owPAiklq/7
pF9XsH4KcAiuvc2M129a/AywNbYZIYOo3NG7prQmAqS4aSq9hkq5E6SmRtdsJJLo
WI5Vn4B3gRUrKBGuT2Hkvy2yEs8r0yY3wxI2FfqRNyfvB6Vm1BxIZOV+gT9BZ3rf
TavEuRDsLddH2hSw+r2GpJ2mWWNH0RM6KVXenD1PSApZN7HFQ7oSjMCmuI3MeCTp
8Hq4/0EqeyWQTmQB8v+JA0y0JmL21qnpUexKc5F3u2igIqmJ0kPgvOnRNFSa8i1r
LJnb+XU6SPVx0pVdP7+6cKRkSyiheWE8H0x8+3yLMBWoQRV5tViIxErDc/bSv9Tn
oiJamoCi2MJS5xL4gM6PsScRReV3fXeUbFcJRLwI3rX2X6XxrqV0hFyBn9PWkH+I
zJwr6AOtyk+bZnvfs2u9V9Zum4xMDAiDahPiSDocn+XbdaJK0tjM3qRaosSR4Zqu
OMH7wQWeQZAFY08SbfDUt7mw+oytvfut2cJgv0JTvjxfqHVi0ZZJgGYdCHiJXhek
NDzqQg6Ijwg1sbSdeluXyR6wtdwYRRVtrVa5vh6Ih9dgE9k1YqcD+pRWA4G4U7pt
6fZ/c2u3bgD+lnIkFOqwgPMOkTIv8Qbfwf6+Hs6bMHAsiu8CdtJWlGkcBVylbBMP
fuERA/oUTEKTjwEom7e8a+V9HDqbkq3f0zA91N9JFtQhr1ppDoIHo5Dq49CdBa8x
l6sVA6sLNfRbPEklzkIzBEgnD++yWBPO/RVDceVIEwHzgti3/0ysWwIUKgszHobp
NGf3D1QPzY/Gel5i+3+TQ1gB1erLI6c9yHW/cPoELFV8RJKTlRS+XZkXBXuaDN1Q
gvZxRit2H8rzdmjlc5Zb6kHrkWvLl8ZlQLbrtwcdpm74qe/mdh8c0UPpSHpSVPrx
Vj2LcjvOA7Asibwc3nqljaYnCvd/Z8otWBKHdBSi9HTmwRLV6b3R3cIPvklhYb3g
SspJLs5xX15o0TeP/vprDKoLvK7Iuw9cU7qSSqI4V0JH2oJcyulPyAnQGNKY6Gj9
3zrXa8fhopSZAku/HmDOChG9mUbVfulUbOC93ZpI/JqQfUcJGUqM8fbHVTrdjAby
rWJP1YpwV3qWaXvBwNMrdWwDy6anxgAtXGED0S2vTnC/XNULQ6o8jCx8ne55o/Ex
WKHYZ7UL39pQwbHLcQ0dinuE+8K6f1HRphoAcFmHpl5vmdmIPHNhu0tvIIt/fUaz
PEkU2iscmb7Mf4niQOVZ1YfTCQxkq+9CJ/f12NYIr0RnY2VGLSGP6BsPavpLSfpz
uzZCD2jwrb/3c0dl8pKsL8Xgryq/Qgk0K2sf5maoFWzlq1dv8jzsoPR0stAdxLzq
HkQX9TqzMes4LciCQj3cv1eL5uKTIh4EZHSJ9VwX5ZFdbiFxKEajPQjTySaO1faN
4yX+uU91AgCJWjguo9HSANVjcmG4xkfra6XS3evSiFvK3G9MpxnUDJiAgyxe1y1o
QsbBH0e9JPAVxN6mtD8y5CVMyei7qMhF/3K/a94+FHO4bts022qEJ+3gxgo09ZrU
eSZQiiawWY3V4isB33ivEhCTVCfJ0hHVPaRKKXyldJjjs9sD5OU9gId2FfXj82y/
W++CdQmt2dzm2Rf9G4Aowsbk8fpr64RhICoacmKytfoyGPYkEepzjizmCSl2S26K
hOp50GkcXJxQHQnHJRMvxGs82tFP7xh7+HVfpAZeVt5RKMGNCPSzM1McQBEtip/b
NlMJx//leL93Z5yIOPSpFmMNLy/03LLPgo3OGxd99JiYJZkmbJ7VPgrJG+UURrfh
/7N3Mr/rJ2grSC3EH9a7D0xYrdlJ36m7MftpCbxvePyPeDoQFcadHoAMKOgXf7Qf
EHGS8wtGrgrzM5AoXGyDZ/2NfD0c9muUUiE45TAK+H01pits23YsE9gB453EQIfU
92p/rWDwPD5QHlGrrKIPedec3d729zTDE8F3T4S/nqFxz0KVq8LnVKGOP9CljC53
RlB1UjNElcRrMW6himP4J8XSElVtZTOSUy8fnoNSG238PbF7wfE9YhpMMWFagIIy
zqw1r4SdDUEwhdttWtA3TWvB+Mc+/CbyFdZDb1N5KntkIIaI3ukxorolYYVin1ff
kPgXCZcRU22vMl+y4jm8a9xb0x4CSEWSfYITHzvO7JhTZfFb02fA19Gr71+Lf+5j
iytbks1R/fFWLoxmsTiWnH2XFv+VcO3FhxrQaofAdp4ZygO4hAAtZqdd2lDFSKDH
DomWdu9LcCmrWvCuAcpgdCH/s+x3my5u8lNylPkJCXqtRR+Ky9pfMav5ln0zSsfP
4OpS6pobcgObweRiHLZUInNT6BXbU9mk169C7U7HVfkWiTE0V3Rp3KoiIVwRI7Ba
MJtYtcH0ShlzSZyAJa6LSwy1oPPBzrNNfxWrgLk/RI/nohzRdaKRTEM4LSD+7huq
Lhdn0xPEdcU3qHmw7UL4X9qT86FTjQgjt8tzT1SXvN4aP8JlqcnzBEStArqOKOER
JrJ7QDGVZPAMFUD3vDbKN0Q/82uo1zjRbU9W/FwMxptXjPVoC3I4+o3eBzvvoRHd
yP7Nj58kA1js8jvBE5U+ZzmIzufNKi3ksIawudvwA8iqKLYfEh3Bq8YDDtytbLVP
acXae8soTuEzweV1as9Fl4CBTiaOa5gZKRbSUAsq3pEtSkfFTbVIDfi+vVCNUpZF
CCDwd5wtF9ydcyrsmtAJOV3hNRA0Z5sN30v9aUkcPzmyN7p6MRYNFpEGAMhypnxD
mwxLAw5VS+E7hxKwS9ZN1nC8E1WldGhRm1roVF8pD2EQem4GrSqFeK07PiCejsY+
gLxpHLIbpyUEp3tNIbe8CBXRc/4wy8FmmoK71g0lEAl8Zt1zeiTizofWTBq5Z6O5
YVtrhddcfhDzQVJDkWVB1u6GWXPLiL+RRNQroVVkzc9Iu+izecihjPDBN4brU4gy
DtiPM1gV4o+DTdH2B+U/ongzFXiSTY+EEpJ0iFBe53sAVaPxKM6aDacwuuUQ3QRt
oUXXPmfnDkeKYuiglLZCDWNB1hpRtqsBHbP835KKbow2bKsNAq0BuyYN1PO+VpPf
gZRgreVKMAtYT6NHvqk+J8LBo8h9SJ+4f2ZAgJEbIYBcGIIffBvy4bM6/B3RDDJp
KK3H704XeMSjqFApirNXfy3IbeeIoN5LDl/5uwQIqvnH0OVN0xzRt40QGW3PWuIo
y3JZCnn0zCZlbgAeqSJtTR1eib4BqwkVd3w/khWM3wVSrKBZGIgPPkI3hj+Xa4zf
ATGl8pai0tXgbrhkuMHOi/643Sc+HCruZegmfC235TcXHR1c5a7iBpBF1p94vyzW
7zcQfkGX0wOaR5VG6y8c7LIOpiOOw3hafpoYo4qkiidvW+XNzGpLnIjMe+mMEJIZ
HhubLIoPTQAS0/Atw81RutvgiIJmw7mqvqC0YraLqZsOuKefh8XKLXSWlinHm0xi
q9zX3Pm1Y7hkTDT1gnwMEFZqAJyTAdes/Bj3jEV3IAttr4UdxIXU5E6UMBOtCpOP
3ePbeL3bGRWtbF3rTHCJaBbGdx0PuErmauC3+3tBmjzNjMnZGvs5d+sWqCXHNgum
lmBH9Y7fydscoVCG/+ra9mZyC2cCB82Tm713RVOhtdv1U5vnnOKiKmF8Hykil3Ff
DzDUoY8XCqJxM81MQjQ6ej7GzEJTq0LXL0eWO3hAu+5KvD02BJYRSPBqd/QDHYV6
/TU/w8eyn9qZ/kPTeM5KP/DuzE8Fm7VBMiMtm8+0OpZYL68sWcDwH46rJbGiCJpv
8q8cQ8KEmO7jtemN4d2qiFDrwh+wLw5JrglBO/+peO1XOSNLqOdCADBRJucpMJjL
qWFtdCvnP1m5kraVKnTzBO9QUbjGvez3cGDhRQymtu9JomKP5xRR5xJOtZkpmDOx
J4siC/tjg+y2c5lNfJV7+IWgqWgcJ9IGiXPDLZUQCM+9994qCa/nGBUZePW9j8s0
O6T95h/POn0y8c62IsUhMMs9PP/YGCgDBfW2lTBADwYChdfa5RHNo0QfTDwswcwo
kXYoUDJNAaX+3lD2uGFMw+sj8IyYpZPc1IBlRgBlYQ1Z+yTMI9BtZ7Cuc6PFw/V7
rxwp5XNI9KQWeAOb0jh5+Y4YldgqDhNyg+GcqlMxF4tYxDOwDXvKyrTf+PxFyNKm
fRoMOh1llqaHlf+SirweH1j+2L+/nl3uWs3CbY09zGLF+DcV7qD+JocRfrkCuQXO
rOpUiVY2lN9Fkx9EPyRmZivJMKxeR9zRE7kEk0QmhTewzt83db52MNUzT0raPIEN
gwefq/BSe5FhaBBtSv5azerJ0M2acFDW6UgGaXY//7OI/Hw864efsXwjDsG/l2mo
qYPFhcSTPkuqe/zAresCPXzzLTIk9mQSXCCaDXp8R8Zx+Afh5jR57PPYiPw5enba
r/TKyd4O4Jj/nAJEvTZ3OJ6SzMZOxrnqgG8O3gVXJ353PjO1svhl1hEb6kFl6wxi
R9zefv2dGMhNxliOytGwNAsKk+lLc4ZOZnM0jeLTiygQXMoTnK/6XE7bKYGxAvLr
opZYLgtTz71LkS2eKtYBItcmakRyPZXp9L5aUjgJUBrlhg68+r2vvwSjAoFcBGT6
19GrGsWmU46579jRVeAfFvaNBxr7YM9wVYZk5zVL1mc7+rjwmSXFUHIzb0oqe+a0
/ZGXawxoEojtqUBYx4aTKFvoivfCPxqwsqA1K23r6Vw7DQnO7lOpOQ4ltHhn6msZ
dv1IZp8K988Z8dVFICpM16/uusEc97xl1v2rM64oQ/ZB3fVmFEwNsfPOJHjFbkpW
UEln9t4vEneZ6o2bO+6doMB70Cpn5S1rAfrHlZonA31zeUoRmTNLfj6zL64MaNxp
rph8lrB6Nh8gywTa15GRzNlOd3TYhYZ6Eg7UgtAlCjOajahMLfK/7EKU6373xwDv
fbohJXIFjlVbzJBPr7WGKsUBHe8cqmy20VzecIegorXmhW6sMVVBO8TV3+mWFtfn
HObxjN+s4BlobTtP7hjPdsneOMsFA3O35pCE4GLYCAJWIHTu53/0Ta5d9FU0rzIu
lzFOFLz6x2MQ19JivHLL8TKioon2KQUZFjTJ7mgjEjKpjD9UxaxK9/2+JWgUqgRl
13yk2XLlqvuBejdsCoEhXfqe/TGI6Ug2blHIQVS0eQTrsYbno/xz5rXlQmgWU/XB
WTeTpvzgXFae8sXfkBC66UPMYs9SaVhHQlttbOETF8uIDLnIpVOVJv6Hk9p2fuik
ueBPppZVEs3y9uNaIE4J+ABLg7MS0K/FgactpFGrb2TT4Dj6owEO23skx0FYu5A2
QuvQugXEbew/F4yRnXKVbQ8+qR4g+etPWmDpiWnyjT/3YyXaHg5ShBXGXzbpwsz3
AKP5NyzmCj6kX5LK0PnaavWtk+QTd3/Di6SLpk68TtykBfLP7SbbfqPjJssYMg2r
H03L0Bn/ksHSsNlrx4qYsiJhNKgMAAPOP5nvV+jcqg2o+8C/48J6XQmkNDlFMIuZ
YHFTIbSBTRpBWpI3sxUXdB7opM+qZk5ys7vnBbX4IxcFk+O7/o1GnMUPpKm2Vi1h
dUaMBxWIgYy1s/SKw78ASTzftZHBgLD4L9H7C9mQCTJAsfZ+uz5O7bw++xebzoWF
slUhl0RYVZ8d2Arqb+/IWk3p34Wl73jsjNw/VAxfbumHoQDcwMXv0MhN/afvN0wj
PH5V4rttA5kCb5O0Mb4Z8CHdWBP4k/JeQJoWaTyUNgNPMESQKIHH8ig0GljqXHTF
KXA/AEsk8yw1Eel6Q2iEqpfKS219UoUbMhLLQo/J6GExNmMW3qTL5VpDk4r9gRcm
r+Hu19vQpjq6LfgaXWQaQwMk+EMs29JXm8dkd9+9l1x0L04+e4MDvmchnkhPTQ78
8sGrvxKxSekv4hyl4zJJIyLrqe5/o8/I+cnjF9IrbbdUylQK9Iztve7HkfP0kIZB
J6KEDsMV8SIRjIE8QmNyY8C129ler5ZtCmOeIZPnQLaKbTY4vujPG0TuaDi95Wu4
ZQN3RjV5Eqikwg8HbABgFlufAQHReiL9Tz0IAyLFwcqz5apHkD+NNEP15kbSYDj6
0FOBz3VykH0EOTm/mkpXQhbjZHcG//XBJ/bMcjjPSvSaG9a+DXiD7dDFwzgeGCoV
4wEhNLMYlA+EnR1xC6mIITgg2+gf+kbKPfHbdXJJM7XD5kFmMDwV7qDTMFulw1Y0
tAtGbJTI/qddyt1w4+SlGSoef3swqYK7v73wOX4HRapTPBWT2GhfVNxCIzIRFKBC
YdHshNykx0kWgsFqA0x77Ph/f/jmVtgRRC+gW1drPVIH57a3SQcRsm77x4Nse+06
KjtnaCmiL5o5bZ1nGLCHccBuYUjGHpGAoNte8BdspA/trwZ3GxYiQbL8zW5nXQHw
zORSh/vQPJ2LC0xHWZsIzH84T3c468t6J+T09AhfSsv2yO1fsF27/r4wjUuGES1M
+SibyxYhRZr5IvH0MwTDsg6Mi0DKsl2X5XNpwpWYMl6U2tU9o+oMAq3GKnnIem6C
gVz1kJlFISdch9M+UlU5edJ4TVgxYc84aG6J2qOqFK7X0LYVCWEU+zMF5TOynMfu
Y/6/cEimTvpUcbraL6VfZ+tf0ZuzHItUfkzTqvNBhv9xPJsTDNQDwTS2wbP61/bz
/Ayts5FThfo3hI6BxABRLH+l3ieC8wwBF2/310d4Z+gdarqOpuA42WOVeoddcgXO
CxqCVEt7dbnEkHm0Ac8lwSTUSPEDbHwfD1xe/NaK0FB8fSRmOQHp3hiHL9hs96Cd
33Mcj9DT21XRNbct5ft413ACNIpf+gzvNhqNoSPjX7lNsPLouVnVEyHSYNh1v8Qd
moB5f3lpNBfHKehB8yKW4HfQ5ex9TWHCliE18yGYaYWskklhxjKvZUAUH3tF9d3V
wQOdkNClAuVB7q/N06eCHq4OOP5H7TP3yg+M8B50ZtVSzve2vqZHo37z+M5FXJEy
95cjRCBoKOQu4lLo6oAp9kYnSlmk+bYRE5DXfGSoheyNRHz4eX0iuHe/mle0z6dn
eQOONeaFXzUIEBE76bF5qU6WK0xJGf4KxUdS+ZOfjzib9AI5UM6NmxxdEHXGkUD5
ad4FmS43u5BdyoWH2pwX/O7sVruaBS2t06CLmop4BwJfMAe73cffIYa5qBZh3geG
EajeS2ILjSAsSLh42XDXpPcvjHCwkdq6kkztd+9fdiH61djGMM5pFvb+DW+L1Xv/
xqXX32z1J5xiqMAYU0oBNGm8RCPGRdAn7dDAjyYMqK4LXesAfs3IhHf5jVgZxOPG
DdfZNznod4rHnZezeC+JWeOT7wwuzYXjeA4HgiEFTgxlIsCqw+Sp/09DNzli2VKH
/bSXqrlDMOxLiXsPZRTJMmYJpLbitcV8ggin0WA01vU+e/UrAnJX/ue/ZevFUbnM
TP7ZNcveAHYOaPJbBFbhWp1JD0fHM24An7I+T6Lp4h65LuVT2gzi0O32NCSAGzyB
ByfWsi4ziUZaqvX9E/91za1Ni0uTT4pRNHmUPdb3Tx6zs3SYtp9dpUnDBZUn0FcB
GEOVrP+KAwwUWnnUScWvcSl2Jel3726Xae+BLiJ4aoHADsZF14FY6auzph5BaHbh
77HwHOpNaO0SJbFxQU3dlnSzydcqhiE7NUyoZ0qosttMNV0d/qJDJotxuisvx9nj
ZzcEhXz+4LEjqWGcML8AcDXPVDRKvgIakn+Y6mHJWIuVRE0dUrX04i6QRO6rVWCF
w10i0hXWDJ/W3QyLvdopl1DKPt7Ot61GSLJ6GATqBwPeVRns/rDLVSc2bnkSJJmS
OWZfUADsZW8lEFdgUzAoDAfvrhIc6BDuaR0EOyx1+ihmULU1zcyNHrABi6xJu/EH
CjYNSa0s8Cy6qxcnyTPqnLB79RJ1iZvn47Wrk8zpo6jqHpV7GfLR2KIISENF1wHE
N/QvJpjjaip1HC2lpzH1ejDvI0VrsM/+CYfYG8CNL/eXV705rlLbbo42en9aLSWe
5yHT3QywD95AYH0rBUA2UfvNQ4fcbM4+Us1T/I4wExjG6cD7xgmK4MD/r5y7fiN9
LMTbkHgsV4U5sk5B6S9NH21Qfwgcw+c0EEt5xBdj0oT3eMwDGuIuDZj5nhx0J7eD
aIKRO68WYwRSm0RHNWwY3CWOkLkXaCODoVWGcYbVL7f6f6WMAiMq67K6gckvK0e8
k+msMZGHwOy5Smf+rrj0bB9JP/Et0idhqZCpw+9n9uXeGLdipJetolTuFBaF3wEG
cXKCDWtBNlI6kVxt6RNg4hqOA46ayhHu9oqxhqGFwR7KhNwq4goQmvDnw4XAmuRF
`pragma protect end_protected
