// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:46 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
F9/PEGFNBbt7OpcSWPHtTlruc1PxkRhYkZpkvHMZdyIM4sOLDq/ko8kxFq98sw5r
X06itCHPKEtDRgnGNxU7iI1J93h+mPY19zjTTOuS4/5v2iD8Usz0QSry3ukWcbkH
08t2935v4yKuEw2G1o6ZHrEVT0pllt5Zv/Ym5hnPl+A=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 9616)
+0tCpxdIo5FlfWA9EFVDV+qD8cXSmUgl4y2t3oE6hMNVvdQFBcyrgoPtfJVIPYXQ
qSGB5VjzMv8R7Pr/8X4ihME7Do+/TZkscXHkV98QxJTLf7oZnN32dVxCUl6ufeVP
UzuzdGoysf8tmPInXm2Y5lpM36cGRnY6JEGdUBak1c6hT+RCi1E2YKXPx1WXI3mv
v06oCck2HixcQdAb8kEvJkPQCUkU1nU6VzMA4+KzxW3uVaSEFCWEcA7JgE/Pxn/F
0jOeg3875bkPrZPZXzmjSzl8fW9CFyvHElcVmVnOZCHYwxjeMAh+BoPTm2uRSgNF
ypnJncGj237M5S5MSRf2SsmWjwmKQVuaILaPSLV+75DrLyhAxYYxS78N11R9cyLZ
GWW6Q4qV2d9BAlPmEVCczfnSHPsrsFThvCHagelnjL2PPypyAqdsTpEpTlR1K0bl
ETFqOEJm/kVGek90tuHh6yX8vDCHMH+238GR+ope8Er84XiKxZYfpcJKiBhpBF0/
8RO5nW+P4CytzbFageW/1b45hoRRoUG8YFlm2+ZUSlKLGJpdUPafl24tKp8dATRT
dXEsMgH0J1KTlreJQGLvaifuYz1NM0y8U6KuDiDzNSoKM54keZJ0HNjzCD9MnIhX
yXXB1xxfepH/dJ5YSiiAU6OzZaTnvXSP1QHj1bVyZdyoANvOd4kiitswXrQCiotW
2tT4ThSD0VacFHlVuwkdbqMbuW/DVNu8/gVHm5duSJSwDSBPBxEPMmLKVbl2PQHk
E3ADg7JQtk72vSB8WAihej/Bjvoe/7X7QFCEQJjS3o3Uq3e+pxv+u3lIx5mH+ING
yrczDgNwMWfFV/Ap/uZDdld5NQjPQIRvYa0gXqaa1pobo+cIf2FbV1dtp3u8JqSR
BBPC91rzwAUj1xXNdbkXFJ4WaDLQn7YAFCUZGI5nbYp3U8KMevtf3FiN+r4kUnK5
iQ8SQZCaf2Cf4Req5WT9jI3Lip6mZ5bQRhKNY/nRsG+LqqpoaM9n7u8qYVktwLYx
ecIttBBG0op+kq5p5KUQtV02wN/JhqUmo7yU8l/708ClV3nnVsAgRh0rr75/KACz
PTxhU4U528lXZjHOXJQ6ZtXNBvyBK9kFhNWN5wKGEGhdxlzbgrKylYA4qqr7Crks
UfUoyavYR9sJQf88gyPrAObGhGBKvPGW3/yRb6vF0E4Kgxl/gEKS+nyqik8k+A9f
MwhxsdefmZk6eA+nZUvt2K1knlGIWShQI0ao5xrUb0/LujbBd1LEulYg5UxmL+vr
Mn4p/VOLUQWXbmCt4OvB/lhLx/Ifu3y2T/3WTuUsniGZxQOqacvN4+yaT5p+I2mM
VIvdSjnzQWfSwjZjkHT0pwUtt5/6u2nsprA5mpoUFYQyiPBnS3cgPKYomMe9Poj5
lIyqPKYhIBK/UPCwYQLtXR9f6A1qgqQXZHA9+WkNYxKiuhtd6sTYttE3b/EC3xvt
/tmaovKWzHDzm9kt5GmnPXGi7bJZVZ3O5EGq3WlxZ6+IRUPF4G5JcsyqPDAuwGWI
RMG39oYYGDmyr3z3FWnuy1ur+iXu1MTEev4OhAogUVCo0UHss3gnndsLI5MnWibc
q3g3cIdJg/DchgBi80orn2S3YwnFd2jyv0bttUbC/QOCLg6dTafjx+bMcWCO54xX
0CGpnrLm+lf6j8XKzNj0HYCDJn1Vbi4Lp3zsSJGWO29nP0tgN996uEtz21iBraIs
K9kSnog0WTVtw5C6P44mKg/Mq1qDveNLPSZ6PH3ipwQ+lFvtYWmbU2op+O3ifavF
4rhgmH87lSpEmbiXePgPBBowQErbNHAr/GBfm6BQseDwmgKCG0fZA6T7yvrZviVP
7zN+mX0QEvn4MC5n8oYUE6Z/E8bCQmgnrrLzVEJd51vEYauPLUkRnYLIVgqWpDA8
y20JBKUvsP0bJPObUOhwzcbwXkCo1EAVJCVGf4eGWSB6c42oG2YXnDuS3KwOdbRr
HOEMEbJKp+/MrpBvHKiwriXWPoPOHKDif67MRFROGlxkMXuZjb31PF5NOQUdPsAb
EToCDF8B0LcGTz6jfiOGATQn+RB4yhh+yrXRltdgj7v4GbYHgdU6TG1wNF7+KTQa
b3xHiuiVea60GW/zmIg0yBnZK1OXFtp4W7dSxAebZt+jCZeHDz+QN9tNBTv9ZkEt
o4y9G1s0lvCQurnJ4yEzHmGSh/II6fvqLA+6r9D0ZP5aNcKCpc5JyLLEnlYDrLkp
Rem0+D36aGOCPlNH/2WQlOlINgGtMKVGDec3PSdKSubazDOEfgTmaBLNaNbVdpgq
LAIS1eGWtRTtdtousx4EtMebarpBGaOiMb5eVon00HtiyURLpay8ebd0Mxbuv9YQ
U45Ckwf4EfwEFee/5G9FEAu+QXlwXQIbGGnc7S+NJz+dgTdXnDCK4Bq8bA9wS1un
EGSpeBWsEZf/zOWiagAdCgCNrlU7erpCdaZwOLZksflArKNEO05zmrmDyP8NpbhQ
jmFFQ1BmIo1i4n2E9bXkrZCFe3wL0A3+x1EnvnFTql7JT+KeFhzWmZkdVGY8zOrI
FEMNr2EDq80/lk3Fwg1vBIokQE5IzbINqrww1O2VRkF50eyuJVhzp9obyFuJg9rF
BLG7eWcHpThulUhIOt9RBsHIfBhBhYHdY6btU3QdP34ktYLodRy4uJKLYWp6LTd1
VldwGvVNdclGWjgWqEam5HqgmURzI0/SkeRQD2kqptEAK0pmXkG89v1Ovo1MxsR+
1x6FQCKWCul/VZM7ZYHTbcq7Dof0FicRfUMj8Uck/2f5RdEc9zXy+8+4VO+L59t4
BPmcnRbPfONIJ1PURboiTuIbysOaFhmvWBuwxkIsifHInX9dyrxa9xQbtJQTKx1C
+28LO2jlVwrfvGWTYrSmDOpJ6ne86QitzhBsO2WqD4GCddu7J0KPBdF01o+oSSPs
hzQkOfs/AbY6QMksX3S6beyqg6q84nB9WyJm/3dSc1OPTtS0YZrLruOy2ph7QYZC
gvezmhWLQdvc1Y8m3aLzm8aRDQDbNe5+GLPN2zFASTiK0ChL3yZzhQA0O6U+FD4F
0g0raWP2YrrCOrTEfEdPox5o9OWv1LK55m6O6YJrEEr6bkpwG+zgYkohohcXgWGR
IIkOtiWGOyclsew8SF4fTmimsholAGxG0lrnEW5noERXgfiFOVt3+GS3RMJQWRYV
mfCWqxlm0KaGhS69dsQjoGW9B6EcTUpnVeXSEgZbgZVEiR5MYqYJQ6nmYBuN/seM
i8wf9DgZ22U2U2gCxIpWjtGH0yHcnMRzal8/CHQE7HyXNdAy7oeweK0SYZXhm4z6
K1vSOb62uJsaUvT93J1mqfyHIgtFPuperkZZQRdDj4+Cml7hL2HPF4NPsnl5NAPi
SkrVu5YsGr2ImNOV3eSI7dLi6moJ+ywFGr60lGjo98rxL5J2v1OQWuQP4jZF72sS
szehQ8nLxtL5H/T7G2hz452Xd6CkF7w4sgCSqsU3R3g+xnRjD+UlkrIJ9OHXOPCW
oS0ZSWIqSUMJZZGnPSzgPcAE0p+66G+D9y14Kre7lr1qA1YILDchVhpYmr+3ghYJ
8/5L+/yUGQ/fcxriMxULZMYBkxeii4UNMJod0UjbByHcxsrj4wobLbWq3tllfh5i
O8H+mgSaav++BA3YbrSjL0WLcViAmQ6PUEJzisfava9YjQoLnWEqpW8x560Dzm1k
6xYU52uhCzBeZkcgnh0Jhgfq8qmlrxP0NWidZF2wweQswEC7FvofsGYE9vKsNRuB
5NQA0X5hHLqB7zqZMZZh0tat+VBOb//d/Ed6IBgxEm42u8OOv0yOJEcPrycRuk+J
f3AgqpoEP8NTM40Hlr3ufuQjAW3qS5azUuAnGTHqA8kWfb56Bn+pElkRCRFU95tW
Hgn/evImkUUM9cdPwvT8aGphCx62YcMEAaPNvol5ajamWO7uWBk1AAt+Gqm0U/Th
Mqokv/684KR4nAnVnv8HMEBdrxI3ByxIo5ZRMBlyI98cPYzHMjUFnOKiK74JO9Qk
/9wJLsqB18FoY0sLOOs4k/f++lvRr+D0eN+c12zm+u+TIiFY2uMl4WWT62bMnSDt
5Al4kgqUDiw+vENBQxiUnbVWQpuFAHXQ/i81w+OgQp6AJYfB2dsnWIKpARI3E8Ev
DJwsrGoZ0r7xjsMLO6v1juMR8mqMpHHZ/ZiucWE26NYNB4E98/27pOEEZifxzCGG
M7imQ5m1vbL4LyUzaDJdcRFJ+0isaxE9MHkSBKhPp/pZcAnA4V90j/wgUTW4xMT4
I94OzjnoomJfsnXE0XThL1RviIUaoSVvXsXHv1lK2GLIiATbnNd24FxjwL2ygDz5
vm4yDF26qiTPklgbrAw6nUlP6AYBhK5hCfURJyrMHsdYlY5zwEAhdAEx4H84wDkN
5KxuhFWGcFKwT1EN0kJDPo0VAl9nwe4p1ESD3p3OCKJ5nesN92vLwQUrwSpg9XBO
ubDaieJuf3Ba0HD4iG2mDYGqLbDeSs+ox3UIK9E0LrELk1dWYuDrICFNy5KARAoV
BYKyMIl7VYlXgYkkEd/HsEVlqpwiMNX9cCfTzqrBJJLhwGbb2gDpWTLIoU6VPNNx
8MPebzrc6nAS/JOTPvRtElKg+Fmwi4RYjf8huftNpsOsc1qj0ad5Y3K8jVbGgb7+
sn5n6DEKslwRno6hkogapsKTbdXabQVft0tww639I5KCMNVbvtJQrIdczUm+30Tq
Af1k1kLQUtT+enGSSsGHm8+Nx+ir6gH6tYfHe8yk+NUfpLXBaC7gpXN4f4nDUYjX
htdNOW8T09mpNublpRgSBc6VtU96q97T0E7eSH0J9wiDqTYDF7nxUBH/Oii97guM
Zlaugtx1PLYxiUjaMEavGxpIdwHf+q6L3a2KaHPIsqJbeDE5OJTEvWGeQIKzdKVn
61jAhoCuzKplafMDmekfq/+klLM669FbFUhLuCEJroguyVKx4EVHa6QWybeegPXn
fpZUANFJ4wA4x186LwtJJFwQ4z/rSNev2aU9MjrLme4Ke+4nQTIpyAsh12kYIFBW
jNR4qahCei9XuSs4lZT3dpHx/NtNa7U1VDUbmAutKkJv0pW9XxSzjvtH0TAXoMGh
Za1jejREeZ8zom36azW1Lw6aJ6YWMR7CDGZXRt1PUKmsf2snaWRFshAttxDIAWSY
B8qvXnhQYYhaHQn1xyCYADDtVsLTt3Di/sOyaOAp6jV0+6P3NCsNan9EUF1j/AyS
MrLFAAS4sao3A4TD8Rw/45BWEUcAg82givEZgNSo9JOUn/xtr/ce3ikqAOMoIrf5
suVWxLWOSvStMuXyXP5ryMgeIUL/UObgC4/wU2hSP7JJ1cse3a4MeX79Z1i8PLPd
2GtLmE1X66i/0RURhNIrZZagVLL9w2cBUV4fpAogw0hrXKTdsybECgtu4siH3+Ql
HaVu8C8mbypdtM6miQ4RQj1+M3MGXciV1JlF2iMW+ErowlTLT5xI1l6XjPLnhwWw
q+8RQlOvRVGMIVw/RwsmJHggooseOVxup9x0sdSDIJJGDiEXxW5Pa21LoRcno1gG
7qJ5DWW9rzcMBbzSUZD5I7wbdqwhknPm1jucOX7CpXUo9f7QyQ99Okih4D0WiGpx
UFTPxMg+bR7JsewRilEkBUzJu46+MsqOr/LtAz9G2fjORCv2Nw7dTSl91F1wWWEY
XSq0FLA2rrnt4QpEnnm/g7hd9HV8sbd445XFdhT1mjoKogZ0jqw/96pUVFHxlF+X
Abjr1rB2nc55uGuFvOHMpza7tsEMuwSlfuzDw6cHigvJR6/Ym/SHC7JXFeYx4vHc
JQ56Gb9P1SbmG64vwT9Xc4DuW31Z4zMgx6lL19Ns8yrkck6+MJBfrMSpenxgO/N6
VNs0IVbG3r+dEukQAmIRTHwAkzpFNyNGcvwdH6YV9t4Nb4aNufltnBTqgiORMrTL
maetHWS3i1Aq079KZcB28tWpvPlNIGPklTsbAxa8jD8CogqWHzdHBrIu9xuEdX5R
iNYxrbtJ/ijj5OGmCuz35cNFp26yxwHpFfqFF6qtP4gHTncHzpuoFBZX6GyeNi5a
0JgTbULXN6jead9O3+tN8gv5xzxlD1GzvicOTG2PmBPtf6c9QsH+KqC9D8wOK177
oBP7okal9S+BJ+8VUhBSe+zSgMvg6ibiOrC1S9MSHt/Al1NqIxId76XCidqfZLEh
QB6nM4RkVsM9FLcqexOMcOjmhuAoa8lGyG1jRyX5Taurbisf30J33uD9KNHOLsS8
ZpTymD4StDe+BNt7TMCsn/jb2KKG4pJfyk0t7JY6QcOcweq6BfHTGBOv1vOosgqy
iO8TLK8q0fpSzsmmzgSpfKRJMfpeEIkvgiIYDdatLJZD0cyuI7USI6ccbFUbrACm
7qhGZXACWj4wRwsMPltc+QPwFT/4NPcUjrQO4mbqYOa3gvKKsxhXl+Coj4xy/p83
K+kFB5D043uLpgF4gnLk93UI4v82i3znJslK9Z5x91ib2lttHHp4UW7IonMsYeG8
G6CqG2MB4GAvxOCZibbsx3uy8Ynxcf8GKrPJC5uZSktIpPfkJQbIuR/8nwa9cNrv
aEyqLrZbwTh9iBVMAJzUc6CW6+aCpXay3NUMzkEg+ysPnCf3FUuAtQMXtG2Decm+
3QCN1GN9dNUtmx+4KZ3KjSMXmEyBLZV6r896kY8enuy92G0+aV2Cf9c3dp7RDxpj
P6ambtiPu3K9I3xFVeS9VGvXJhvM9AfAVP7iB1S+6sR/QQABBY98etAOL9j1BTug
/nyqHQENYEskS3PH9baNT4z4Sq1eGEyprzKv8xatBpAKq2aNhKqkpiFzMQoWE313
HhRv5Oy1Y3s/tpZgdEen54SUpSiJWHxp/zwwk1cwjS2ZzrsfZuYbxoSQ9/HVR7Yb
ZsWoXM1eETOWbF4k9s2jqE3gkJ0SdWOAP8XuUvPT0XRPh4hCLw4Q/rGKxwrYZ2iQ
s5z7kiSluSs97ykD7qsZXavAu7uZ0VmFr2/OFkfoqbN6LH1hRw5LlGyi+9HemnQY
a/hDmzUebiZCTNzTMcKs1IEdIa8gXzr7O6QCy09S8HskZIZyaDit8OHGr+du6VEl
Ijhbgg3NRHQP5i1/B378Vxw88XrpOnFDEMGZ6hjJmVvbA9OlbAfWNPuCynRINJwY
Jrh1gjz6bGKONPXej2L+YAfnDj3UBMUS8H3fjoQ4xdOLWUYyBSKjalmxoMA+UVrD
V0CMm1Wnp+iCrxEbNbXW4conk1Y2IMMQDg92rl37727EmIKkezDD2Y85B5DqOFLX
COQahbHpmLHHzpoeDNNiF17Fto7X2Y1cZJx56UxBmlchnF5sB4AxF4TfFUIccLG1
ub2G3J58Y90w5ys2Pb5pdpsgmLKmsSrReyinAfFhZ1rYQhF+SJ4AtSKszMt2X1bG
Zno9WI27QQ045Ue3Sx9hdxV+VQVdGEP9nqjWipfFNncxUaZLFt0haLdEWtsYXnSn
pFrHxKSwFnMTdltoULwRYhqTr3LosKI91HXV9//1ecO0sfpE3PYQez4KMS3Z/A5D
rYRuaSHOxuyAdL30DFasurWVHspPMAyP0+v9uIBQIBBF0p5r1+vnzSzdq03H7QEO
0nSZQfRmO/ciCJAnYreIBhvolZRtjxzBJ/O82Yi6M2k5pBW3h/d1saJdjNMA/h2F
EKN9Sb2N1DAN3mgNsTafIXau61D+rdRfhRtOWGOOo0dddmjpziu//8oAlPy6vuHi
ULNzpEPuHfwKLCXmH0n20zl4KgxnNIrmdc9d+e3Rc2JDYKBbQWEPaqC1ZlDLtIS3
IEv18l4dkJ+4Nlsvk/5CLDQ2ivz1BtXv1eVGIsUs/YCEPmQzptKXbyi6qzk34J1D
Zm0LVTieZt0qOVlUbiLvPRFa1cY3QwjYZ37CxPcehmQIkIPecsaky3bi3XL+SfcE
9ZuUetV8hTFxFsNjRlzZSozzoDNzNzjmwW76wV1t/EhIgQfHnsTCBzYqxhvrtcBK
G0WVJ6PPDjKcKNDz9+x7dg3BeqJfyZ6ybUtc4DdlSDe9BfptDalqAyD0ZGMWCFFP
mCCOKGFSBihQCd2WJMboljGFVIFJvrVkjALWEEGMxyjZ+qB7MjeDqxtYJ5v8Kkd8
ehhCFiGWcAa9LM2T2xbW/fmms3h4D8sWOxPdge+r4qEM9oQY+y2dIxKjtTzpQKcs
kBoBXUCKj8/2yUGwPcrpNf5k+sfmkwjC++ZnFhLpqv3P/oA8NkUZG9sTsruX2a9i
hVJe/y/OERY5bBZkA0NRnQggrzPc+X6XfyAOeU2D7nWEZ4qs9YF+nhqrzIXcdlU4
FiY7KoqN9gLMvcGEiQ04rqSf0BXbTrwKgJJnEkfJeARWcLuO/nucOEvmxFN9vfzN
uro8xJi+11XP/ITDEuuSiI/ry/6kC8hlnVEa4EH3SAYbK2+mHs3ZQdgrwgw/AmgD
WVfWGUCRAbXDna7B83KbPYsvld41DCGWtRlo9+1JctovpBEGy7f9fOsTZVE5TOfT
hY5gA3KFETAzgNdRIEcwwZvFskBySJTuBETLPf01m9u5RiXSFTqLm4yrrGudk+6j
Ilur45HfTGvt0GY3Ihs21vj1XkB4FSr1AJ1S/eWZS8fELhQL89yn0IZ0G3rBgFZl
OHsJwIedDY+c27WBeTm7s/MEnADRuQihefrh4Ki15LEQzFTaZX4Vem1mSXd+HheQ
Vt1R3bVabed3uoT5gvH8X2pDeM/Ijo67VTg52zl+/KtPJpkmHFhA6K//899q76cb
PmH2FqxqXn0/qGxdaWceLclBrdtphSRuKXWZ/OtnJauZ925rBpClytLyE24JBcse
b5q5buDZ4nUAWV2VUQCdNOMD0N97kB3Gv2SyNMWGhBjpzhRfhQHlRxrL5CH3lw5R
orYNcy07CrQ4qOHKXdoYt7hvOj7zsY7d+V0XrDkhv+O9CoSyH3Di+A/+/QxTXuiT
pqjt0GKbpxtEs9O8hcLbrs7uWHAEfNRTbA9InWDIg9cQLT+m1kZ8lqPvD2MkNkY8
zo+oWgHGkUGrsxqvScwj551Zmsf+RVVhQwfFHiWRariE2pGWj6bI7GboPoQIZDYp
j+XD3wWD4cQqP4GvVD73Z5zo8kPzWyhqQ+yMIAfeT4vfX3RKb3A9W4yV2FMr8Ypx
ZjoYnmjbePtTxiPO7vAND+0lFlS0Tg2KmvtYud/lheSEf3HvGVhAIrqKU85qx7WV
0Vv2GOmJyjUtf6w2w0fFgDqvA/Rs5cMEFEtaDUwzEX3lJzlpclpUlurM0K47r/Sf
K4cENHxZUvnctQsKnOgwPAPsA0XcEtRuKD7YwVT0wZZ28Pc1qxOJCxuUXkyao9cd
7k1WUsf1Ow/wfjJXZWibFsle5JIeTbB4uVdsHKgiv212kWXqVLpNBKbCNJdbVXrj
0UZD56LRl6Aw2jn7ntLELDoc4W390/7Ih1/LKyYDkq6PLWdZC6lT4GUqvXLSywJz
KFKUB5TyC4fyykIXEWCBi29vWbxl/nPSa1ielLozHQI2lojISjXMaat1Jtws+Hxp
y4MS6Kk944BPQMg05Do+Dpp93SGJuvrRNcdVvsyg3JBSJfAF6pKyBt2XhSimJflH
hPThC/YLp7e+sLEY2x/8J6nlAIAyLh0/Y9qhnrjZRpQ6wUe+NCwxnpXu3X9kGlA9
vzl1bfmD7VFTEOFyBtI0oPA0eC5y4s9PLPc6t5JQYsQa3Jn/Mwcc8O2v6BPYOSEu
ESE9SSYCUB1kx6RbY+soUex1pBnNor6TVLCH2m2EOU7gIVA9X3x8Hgap8tRq2uVK
x9Gi6QOgNdPUfm80yu4j2jYo93EuePnkcR3Rb1FuC+QQOVVVFrqd2jHhQUlg6mRa
yirLc/YED72jtmI1Iv6IiTqWHLqjMLtd0u1izSQAmERKxbrO/MpH/8p1W+sF26gj
77M47bxTty57tVoO8mLWO0Tu9vL2GROdyCojJcXYGJlCtfWK/7FZOoKMz2UDzq5k
p4crOeMnd4IiHlK2YuJ1Sx842mdDRqgIMvJ3pnr/qFtcs9SpPNoMwqXMGAhW5yIj
X6XrD5bIF//yfOpkA0ahLLnLN1TyhR9MrwahyQTKgA1VKehbCm+eN2hf6q4IXWq0
Cv7UHyVWeyqr4QBA9cOuokv5b0bIWekxk/z1ic7Xdq1ryecespP/b5tQyXgOa7cA
Tv7Eetkc+OoNR3SaDkXWDCeskkJliFfsLgb6nVcKlWBFEQjmlbtg+iZbDt/4zJsx
NcJYUMdT9q/qegDn5xmwqIrHrBSdGLc4hKMKkezsNKmMj1obTe3wppPfoD+ZZnjd
0S/rPqmW6YGwvfyhPRv2Y7QY1DRY9bUbH1ZXQu+zfv2oPlUy6Ae4PGAlw8qhPtlw
ojYYdwh8enuCV5T7AtPPaI1O3arXeZtcpg5dm0y2RdxC9fH6Sp8EI9OqtZ3RhWBx
hBLh1s5+ZJf0k9cMuROIoLxmooJG1skdjMN4PF6ioWKyAFy9Irtq2Kna255viXX6
QtbN6SeJadXetI45SVeG8w+9E5WpHkZlCW0Tks+wRMtWH0zWp64twGnpgEBvSxuj
c290aZdW2vlEVjTIqdyDFeWP11bcSRqpozCoTYEdx7xuSwp3gu0y+fZ/+/oQlZpa
40yE+Mn47YJAVOZGYXm+ScGvzlxpMRWPCoT7iPWLexNHkf1mSPixXzolOJvVmHno
A/xxFPfFG+6/sWDT2y+rJuQKYQ2QAjyv75vS78CtU9B8MtHPVQbeo5xcgGlpQkcL
JdVIF5wGizj16y/zjzXuuG+EmzhhzsFG9ZAl6V5tuTaoOqrir66jYHxsbVSBtLLc
q4O5DoI92UkZERIJViAiru9eaYhNFJi247NqGpTBCUnv4Ac2Aa8ziqrMye+GWkLG
9ZzW3AgZeUDYjVQ3bRlYhVR0y0g6Z+j96u/m2CmsrUX/JMme1DtRkT0OvuvIpwaz
61cN1GqjUW9NWHhIIuUJKZPrfEkCbjQvQBaLuUckDBGHoTKqB1OqimVvTlzk7GIG
gpXdHHpwe0iJ0Lh21dJPnkmVL6KWODR/VQajIEhQ/wfTHe1aTpjtm72f/FbH+h5i
VLPIapaXbpXf824AxDRQ6zZGv4CYl/vUXFLj79glwsFV7Xg9+usjuCRnKeQSkDK1
61ZGF39d7KFkMTOE+kCvpmahJO1cYD30O3E2SXaQy9C1wysK+Gf3LNcYV2PuJ2JA
PHr3z5uC1LU4OeKOd36mN9liurBn3astcxg6LWLLF2SSRXilzVJACiXG34f5Fju4
/8E7SS4kYiFvuKBHv6e5/1BnlWJcFz3e/Q/0o7pePgiYF0uJDmnj1wn8Clk8LK7b
MPjRI9cq2oHIVoVmZXjWJKrVHRIuANpPs4dXetksDIpjTA9rKSyiVupHPPtNL9fy
Se+bYSVCwbPn7SP12tgzW6zG75crCKh71IBm3rOhSwSABlz/yneP/t7sIk1yz0l0
BQ71QQICzjy13sgzDByq3ENIOC+CbrpY8M6Fp0nx508qK96nYrbz4Iy42eKDwGr0
RdEn8yKNW7y087ORjlJhHxZkdaj+JcmHfIbJvn7wPhCypRKmOt1LOcAEQ//GggnH
ma4MFgW0J22MRncpMOzloUe7FW0chHYuuLlyU/uarxUjrKMR7VNqAjXRVcFM/46e
inBgFRheG2Kz+yEYZqcgrRFCr0m7JydYTRyo7L/M7jGNZdBkcRnIP8zQ6RQ8cVRm
KZkbz1Y7lcVZvD3u2zq2v565/PGyqBAmOff2HgyCMMNEIboTv+gu2u/Q9OXfXqk+
Cscb+eyTVmQXciHPSRtT0exweM8S7BoDdlt11AurZZAmjYREit6vSdFJcFpS1wNb
YNcsTkJThN0bhvcadJwjIoHqdLbvC3/ZOhYLKZqBzzV9Or5ZYt1WKoyOO07Tyznu
QVtOnqmqh6xbAWlzP4S7fMTlLFGum06tK7pfUMP+IT3gg8Rk8WyHkqTojwQDaXda
WyOmn3poHwtM5G+RYRks8cYw8TVZImrLXrF1IE3e85QSabwexT2lR4hI7wwy1tL7
hHUO5ECZlIb/dwZOii0yXUkZnhEt6d2ebqJWbQbqbtaVEDHdOLHAvbaYZ+Da4oN7
VV1WSdeRuYRxBHKrV50PWjQee/sF9x8nKA0KQfh4rYAEOTzj74+hIIyDbr4ug2Fq
LDYC3kBgAU5fJICnF40wGmWm6KrLnagYBUOr53I76o5l3KTVXzFsoexb/pnQ6byY
8MdQ4suJ2dE5BEgEkVzqezaROzi8+aSw7uwiFLJp0pxoh3DBbzSnT/FV0QLNM4Wb
ALDi3b5B2gew4xneoNG67q579wTIs0QRxRUAln/t1uy19U1hsRJ6QC9pzyqIUl77
2fnERee109+AArbYTalC77/bX9MdFR8fhBjxC4J6wEEvo/X/XS3pmE/e4oekAYqH
nlRfmrh+1v/jczM2tlbW+d3S++94hKN+r60HoU8B62x8Wehn5qlZ0CeXNWZZLX6h
MNhjdSCEMP/YtsNVO/SAbnm6REnqu1hD1a22oZLQatGm78HzroJ1A2a6o4HZQA6J
WgBwjYmf5kmQQiToeKV52A0nflXjce36BhxPTp+LjqQiqZJ8+b+ptsjkPBD8hlPu
fN2Y9pH7t1EmgxYHAxADT+ZvEavupB4D3/BQBpz8j7IsiVBAe3kie+68lqWUR10P
uHI9KT5k48GKKfH//FbJGJoCIjtlYqlQWae+JJMhe4EA6ZDHMWBnVMsyB2zE8k1s
zQo8e9H6j1TP3xnQTUbOc8YI2KICJJP/aivhaz1ilTD2QlcJ7M1aOj4Cx34iAbjf
QvpFI9g+dXI6ph8dcU0CmQ==
`pragma protect end_protected
