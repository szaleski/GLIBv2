// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:59 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
fn1ysKZ12fttKx4lpWXQBOMvH6rt9LWfwNCYrUsBh+xtSK8V8s15K8hG9mXy3sEh
8WWw6IquferQuT+qB7EYBCWX1c7zOItwdBYVAGlbTG7TLgx/5mSAyae6a6zNW1aF
9SmQkG/IQTJzrV5lJZE3HYz0IU4UV5/fVH3DLsM1S5Y=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 21984)
Czr9bWcwQ6u5LmBYVBw5KDNuZDStreGk7TgTkVprpW55H5HGblnyvL2PoutOk2d3
WkCDk+8eq6M2W6CF9JrSJ8n0nRW41iYofzJD9qR/h9muekOISiWnG9P4YzrHeMgc
Dc3X2eVSUuMRpYKM9EXJiJxIzJCmNyDNoyJkKCveTjc/WHSesh92cDAAxuocPFKt
SITNbgkPSH79QBRwQkFKz8tjbIQceq/fuCaFh/sHWF8zNwyrCiSUnUfZp9XXSE5U
zwOzqQXo1zYada8vAFt/ya2pXARfx4Tk01bM2vYW66vC8bavKZw9XoguBa85zO3C
83jIWfRN40PvOyHCAREBYVYtyjZFQR07tIbdU9cUMj7CQ+VUCTIk/2uMZpouqnMR
vHOhiyaSqnNCHaarh7c8KSvRLiXVeh+/T3cL+bZTrZZsHIuE6U8lBHb1RELGMNMb
93tQ+ksC4BNrAHkhRhyB7tphPqYSR3O6aL9ZF90N6r9mBQwnKK7+P4QOHWPtZYIU
5VbPFsBxeDEWn89rWF2vDJE0up0Dax1noJz+4y5YXV0kQiJr8p8oc6lGdX3Q+Te5
UZn1XReIJGhJpDqVLHWA+PG7yoZSOm3I/dfE4WlxnFaBA4gWsoFJwSMtqFbFmpRB
jYQ4dRSt0WQtdcEpWZsK1FKtgksIbmUsYhKldt5zzbz7fhXlWAEppUN20caVmqdX
4Vr4Z0SPBpaoT8qoUbvQHtWl+PXmvWi+MA8vmbBrmELqgsk/RgRW35Qg9cXFlD33
5I1QWWPxvysencfXFsJqwj+moMJ0sHpTfHDJ4PJpgn7t0Q7y/KmegKXCZ2aEbNIb
Wr9OPyzx8JF89Il9KKGfVujt4nhUL9qSKxe7rsdRY3KSCD7Fo/9IYFsVxCp4GWT0
3ROyzK11E7BZ0V1kfcyiRMdmvphH2donWe0m1v3XzoxHLzvHbGseZFWyJMnX9/DG
Z9Sq3g2voASRb2oBkkkVYt1bfQwNH3aGSZsWJlv2ke9B70shGBqOsPi4bEaEqx5Z
gTQ6et+G1gkmcOsEe5Sgkc5p+sLp1rUA/RHfwzouQEJEAYqJE8xZJVSxL8P7IyG1
ThP0s8d+eG30OC+MloiVbKkxGP0VGfAIlbolBWAC92MRocoUWUlOCAbbUEIBe7h9
LcS+dWxatKPvUp9TUQmJGYbazdM6dnDlkjM6oHnADRKh16u9+uWb0I+csEeQrGm8
h26fXdB6sKJ8e2p2gMgi6LafKTXpTtldvljT8iZJbvcfjdHjgb7HAA6pOcvACI95
DJheufEnyEN0SgRstqUoVz1Wez99wlPzqfriov5Y0hZh/oeQmQ6R/RJGrdAvxLbM
kQia+Gc4AMn7FNmGuBpzUAwLUWiJWbLPnWXNldrBNxVgpG9emeC53PBvP1QoNNbd
zt+OfFBCxBEAgn12w3Se1D1wStNewicOEaBCi/NYuDnNvicu7+VG+cPot0Tcqg7B
BmBMJOT0UkwjH7QcBOHlLsREDIEe28n9RvTWToRHNmiDSGHGk7+K7/03nIaWFZ0X
2Um7fe/lhELVLJY5HHEb1Vn5sB1oAr7xlNgfZHhKBA6RqCDi5qzh1xKki0dyisGH
4qUJZ9ONVgO0pUfwR4m7mQt+SR5V0T2Z/jvkO9061R8/Chfldl+q8OM9foLKqJ9O
5bN6y2E2qxCwcMG12DRvTmVOU1ucv1//c4JOUeOofZt1neSLI9FblovAuIaDGwtA
bstb+Cp4hpIgSARSoJxSWNCTGhLcgab1oKHcsNAr1uIX6kyOlcUCcNInArSaLd8X
UpHVr4JxW6Auhv3gc/9drD01G1HaKc496yU6vhSABngsC56xskVCzPZvZcQXkczp
3ehD1RMTcEMfMpulAYxixeUltjVeLaHIkxChsvABdI1j1zlPMud8/RwrsMyNEWkH
UFyYo7MptxuiROBjcTNDmJ3VhQR2+clp9PEJ+gqXz4Tu2vaPFfcFcgJAUrXxkBse
SX2ltwjnueRLQree5YOIu9eNXKS5vK10rOQ/fsFsFT7gs/8FEofBQiVQjhkpGy/S
qeDUdf0d+rBvzYq7fJ6jXdYUEVSp5MqDb0z2hA8drRtM8guFo2Hml3ieNu8jJ2wR
z/1yeNGZo26Uyzocu3tPNwhBqpzATY0njftfBzPzv0P1l3+BnX+s0j3M1ifsSZyW
Lm4ywT9w9qHPzh+9tQ9P0YsEQTPpX9jwux1RwAuaeROvYGRSaIGdORzvftiNGakg
S4acMqH79cY96ReRh5wpFIRAriAY54qFXvUyqNuA/V9L8WV+WkS+ssL4uyosqonc
GU0ScQcOmE1kdVB5yNlrjvE96J0YQ+H9ZYXyvNhC9PG3gKbew/iAqkY/ygKr5Fa+
ZxcQezvaYmKYiTl4w6rjs1osfLQGhfs+ZhNXum1rLmcz0rJ44VoHqtm0afU2BJa8
qihVLgiGxSeFzoV86WFe8+/lBDPGQVFSogJKI2xxDd5GJaX+g2JyTGWxLMhCWYxd
vjmeq31iRyTzB/GZSXKaXoIuGz60cHgLCgRdLFhGsc5oxiGpH7L0k3fwp/XPNVso
km/T022lvope+wL2H6QkAa87LMkAvvpJCUBZZLDFL+UUxmE/RrbyPLJm1hiaYPaC
IcSCOin0f+wEUWPhygIEHCr/oo4CsxZGA6T86R/q42oc6/9ZS4wfAF0XBgen9Q60
BcU7Gjtb/XqMtk2/nR470XT8C4Nf/1mxT2Hye1AVrEUN3GiopZlzNpKaPGmMBx+n
o/BfW6KvwCcpiQOhsJ5f1/BWf9Rfw6ucYDujrDLPtoWGOX1VPQsaE0/fMs0W3PzO
smsTHIXSaHKbZAC9U84Lm/urSW3hHLXs6L4+cr7eiYYcmHQfDHVs97dloR7laQ8U
5KCW2qDTjEfHal3QFuAZaPU1Ca//aEaYO5nNO78qNGUNdJzP49B+ntK5xSc6B+8d
PJt/haxF43B+kknFql4EYNpPB/ax5deJbmYjy9qQHHeMgCJbXtACVGbEmm2TGXCk
ygcInDfmsKnYXK/SNY72lD7WF0/UWjAzq4seLF0qk9oCA3YOX81tJvpvVEvjfLbu
BkPZweP7vCh3cHemBnJ1IbOPD/+E9MrqXMzpFqu8cLYz8x6MbXw43HbY3psX3w5a
Cl6DJ8oBBnQwMsUed1luNpYKJGTiRrCDuI4J3zHsIPGPPObXSKHwlIHIKUUk2IPM
oimlfuP+c/Lo9Bb6UjcXhh24RCnJdDTUjd5MWvh6xySWC834ozb78mt/bYHc69YT
8xU4TB2PupXq0BwjqO4cElglQkS9PgD5iFNuXp3lENxACL36Na5m364PjEKYul8H
USfivT3TjIFbHkZzWVPyBY5yTRwdrTGlEeP7oCbl/yLNg2HE1rv2PU+8G5BFNYE0
ISQxJlBSKtmvKjYgHNIdvyqtN1rfUbhH54KZKQyWRVflvZy2RAiAeyObBl6J9FNL
Ooz51SgzLRLD6Ioj2EB5fCHO/JA3ChhZIVW+iMb56lmlUDXCimctg2Y4yfFy8IHf
P3j3FJvRpMQvmFSIvrPIP1Y6pMjhbZxavBeTmpPkOl7XZWsSY9FuQxq99L+Em8Wo
MwStXUqME5CsGTshYimal7IQKIxdWK5+1Y5cExviDivAvMOqCIF+htyoQfy2EIU8
k56xXVT/UgUNE1ogx8MGV4tCT/cIW8WPlDvlZgN1dCBQBH/NIqw0duBL9Yxn3l7z
dyZbEQFUiBp8Z4WL4/SbZNwyKEf4G0bunHAuY+op43xxNMH70XiIJwQXCbYtXOfb
l9KesOFKxrsByvqJUISeqwxENf4ffjFLSKWNpfNuZYBIXIYYwtv3XmqSozXuP9Bs
LdVVtanGJDTpS4WQX9NhgQCBmj8e2AUscme9l54YnE4pfRl0ME6jcjLwKY9ED4VB
gqe+DeLjV2SgqWF+qRjBuwE2RvDZXP0kt0IlJqOz085zUpQDOrSr1sYmWJjNOHQ5
tMWt+SKMaiIswP3tjUUm4kiikWBP03MEeCi+HmZ5A5mLcTkq7pPEIZ4c1daoRRJT
p1A+OeZgW5J4I7KwZM5Cn/w2GRaMX1B9V03uHV6SRoiuOr3Kb9uu4ijVOQYTvn6c
mB9CKTC5HsRRRBk5fhQaYb9L4muxk0cBtAWFEUuBn1ZVphDI4t9yGtyB/kd6OlYk
Scai9a0xL8b2IaOCmDUraRyxZq+bahIUsabDFI+9EMweX4kf4h2o8qy0rPAgdXDP
tRrcrPthUrAQO2BzEyahiZz0hTxg8zlzqOHfwLYc0gR/EVihiNORSWK8QdGpbkTd
mfZgzLOjwxqaaI5fR6d5Al6/rJoeUQT0lwOtS3GSO14QeeQQ8le8AFhn+oWZSsPg
UKLXQk/2MrxcfNNp1GaCREQj2RX9gbG67fa7+qSezYVASB0zP6y2v+d9zmbQKuap
QzyGJ2BgULNqE8uShAv6kYstL7Vva9c16NCvtKoQvgpjNoURt+Rj2NINf5eoUM9x
CVQnzD1Lj2ze5lt4tXQwQuvYd4YqvjA6cOUIfoMYPoH1x4SEcCsWc7H1/h3ObQnt
vm6Qqd77HzJF3V0kk34LQ7KH3LasMbFUnKZ8bGrESHxwFu+ZaYVgZQvdeMW54AWk
tvx++wltE/VIIzVc8B+UWPJYoGhoNC4YfWVFqfhe9Qh/FaiffWzMKhFqhHW+J21n
B7VtrPKrAixTlCzj73WSDO7NJv86M+kkvy8MoFj+rF1o8F9CJdWAL/dQagoLYpap
TTRKUlYRdUgtgzAVTjhcq7wX19MpdDw9ZBqbND7EWSRzvRlZj3wEgIy8LyUz2Wjh
5pOQLcT1BfRiesYibzG86vKOnsv3ZX79rwKYlfdZERFyoFUrgurXjFWiuGuvP6pc
w/TbFUP2fdygxKvVK80Jm29MmhXKkRdDThtTAEE0nNREXHj3n2mVDrDOZgCaCYdg
qBEIFM4TmKRezqUz2yyE84pVLx3gYsyXCLS/+eoHSe0OsCOLYPmNIq7W735BZPfN
J7m7a5UD99DG6I4b1n2ByD73MTJiMHZ67OueM8N8mJoCZjc0b71ft0aTvAWIWOMU
qKmm3C+cuAAgBu1xKDveH5iqO1HMrCzQHkgDIXo97Ct0qJn1gLjPQ8pkSyOjvKWm
eXgWb15cZXqt8u6qEz58d990YQM5Bqo/vDSRNhERoDmaHh+9p3Qbi1wn5qGNtApE
sT4Tk0rG3DSyCe3cBWgzZJ29xP/E2XN5cjExehwRxR5qvXCju84mAj7fprmW4HXW
cgXB9THdsu5wmuV1Qs7/Kegcxxb0KeliNYLPWZvbQOdsCGldlX5qm8ItzhQrNDhc
3xS0Qnp4EH6nEIOvFZve89aLdQXeuX5908/iFw7VrJEXQoISL8uBWFyeHGLp48+x
p7RBzjt1qOuh0X5lYCyzAppX3MrFsFRWw3H/LkfkS2xIVXMvihuIXndbOQviZwaB
crOj5bs09EAU7um5VwQd2aLDo1y3w8knWarbx/8GJyUiz0/eg4Cjh1ipPa37movh
rcGB8rQk5EZzyEk7mrPhzmWJnooEnaifsEV7h9Uvf1xBXZy0EH5ryd+z5JK8rche
sFLbbDCAhXprIBHI5WgY5WH2n074TuyST9x98+B30WFk+alGDtHTE/7VKjJjnwS3
1Vm54JGo221Ewsza0/wl0l1KWh1GYvrS7nouBkeE2H2MdkDoQpoEspo7UI+qELua
8nFjYTyfq8txDip5XkRJqJArAlXUH9Vv5lQIGHrI62UMiyber9CBHZzUJAM+Ytx5
ACZziTIa0tWKIwQVBEKak4JieaxHfS8Mpf2PTCmwUHBPeelbzGC2l0UhdazspcnI
ycG/ZD343M6RTgRipShLPYpvScqJWD7nwxbpMZbW+VyR2zs9SxwdRtaYw2ijzpZG
70LjJUaS+WGeuBP1mCm41tR8nHLkGpgVxJ41VzhNMu1Qi+m949XGPIwe8r1qLc9v
q5zm1ZDScEcWUk0qs+qJhYsXnzVpU3Qjq1MrPfuotYOd/ejPN7sjwDjrK2DOSOTa
1NxQuB4Tk1btxKFelu8qc8NxifX23N94Og0qiasJOb9BdolBWii4jpxOFLkhwaKA
1HyZborVXXuOIWBQ9NaZXiDWld3YEjT/NfWM/KKgF/THVz4twOUuWaoaxrcOwBqH
mhC2MN7E8GQ0s+WC9mmxxVyr7iD9eWVgSzpeqeh3wzG9Xf9P4eQBPRjkIR6jqRlr
Nj0Ce5Mqq3tLhO1an9Lr63lzGoM2KbhSEw6mSzbzZ3Eg8r/cYR0A5FcUkzH0JZUL
RmJAgjL/MUPz+vTWQkNDdEr/rMJjeZxul+GRQCMQCOn5d+vSqSqC7bfgj2nf+gVr
sQqN0PSLI2TlGJ5qeu5/f9+JdgAJIRB9sDO+pS5ZLqDDjjoQdddX075aZaZpS3TW
UHQsBfaXp/UVt9FV6/oMmnIEVtUbFNkaFkaGZG14EewM6Gq9M4iMW87GpXPb6/8/
v/JTrKjbpOV4scvfBpjR3CK1NBr88IGl5m5noewj6te4xQFG2fPVfFoaANwhSWBf
JyfW+m1hGFFGSy1whcWBUt6xLOvvJYCDEI+5tPiriLKqItsy0+eAwZ43yRWRUYVq
9Ufi3XrfA5Z1Csrz8bGw6Kh9KoqJ7b4uOVURT18y84QThXVC/bnh/OLUQW0SDTX1
fzoBPT+5PhkOCyfygBtsZaSB6lmyTdLrIvvxZAQWvU2rHLwH8/Xc9Mh4ev7pp6vS
yJhtkfBvPYditDemdRSxXswRvvrzsZdztattYYqQPcS5qVUSxSAGrUb8w0AoQBKV
KruJ1tyjffxyq9ElgYVzsrAnrDdchMv46uKlqPxJUplNAAva52RbGeuPC21VYDwm
HdGNJtkvaeeVtaZ50wcnCO4Pqkoklw4bDw/uSVxp14NW4JEpvONICoIHh6BjxxIU
DqzzV5prbcWnnWCV4C9Kh37KvvQurovljuYqsI/u/aJljjPpsP0lkZTSHKmMTZB+
eGDjVv4AsDm3dzO33LguDfBI6h2Y8u/cnXIcZaEsP5xyF3cOjuVJRshpzdvqyx15
xSG3oGrf/EBUcTi5ckhRgY9BYIh9jy2BWzPB7Xgfxj1m5wbCKXQ6X7qnYWGBtWQD
U5ZY2LN2s+DkqkgmE8/ykmhaGZizRY4lZrGrB1Hnq0TQvSFsUmIkSEagPfjBxY7L
91jLfwlQSLLnReGqQnIHyfziE/aGX03dJx/lOYgmHHa2M01tJIE7iM0MlNxY0fqx
opR3N3KnNWLQDD/PA2xTftr6s9+eg8X+KCoNfP6VRfwfha0CQKmgrhtygar9svvM
ymFCQkoHMMKMkrQjLE9NwQdhNS8OtfSN9KCPyhcvArl9Ap2YGZ4tvnWZT1cFL9OB
GjvsKwsv23ZhHThBDxTzYeuDmpZZLF57FnBof+IMcc7gjInLH6TsMfjZ91b63tKg
VLNNDznb5iMfu0FcCBp/93QxWVKjwq0znecWgOweAK+ypYibD1V4nyrf8cbXcFG/
sWi/isYkxD6Y2C1DUUul0Xt0s6HEllG5Z8sGXqehEIcaSTEE0kj2A8Po9GTPzM8l
CoBug3qC5tw3e0SYTwRfQ9sFofs/wVCmW1QqY6ZqdHbyAJgALHcqfbvJyrFgTssK
fm5rPjxloWXvHmlXelTj9BCsdFi+kCJ1KKJpb1/pRJIIMSPPc1TOKGZdYyB8FCPK
Mdn8wXRdqKEFZEmbMNEvWvL7gDYZwmXCrq3OluKH4M05CGEiuJpQF6AvhBKrTr2a
HKUCkXyzzDLFZPbntZHKHx50eHuTSpBe1Qc914JLjM0tirlORvL9fmfPWHfhZilt
NDn1+ybDEWL1PyAWCpqsFnDW98cl/UKwRw6oGfK3Vt3zaX4ACW5gNhglPOZDagc1
gDD9G0gJ0FDUJjUkRPNR2It+5GpYi6x5gh47n4tZla7eHMy0Mc77I1G8d7/s3hvv
TgtWzZllSwhJwqZPzfzdxUad7ZzSk/UEi7pLrw4eLrD6wjPOhgr3xEqo3R4NoSH9
ZpCxfNlnz4CI5QOUGJcqWeUGyazJE/pCn18Lk0iHN95dxs3e4U74i0h5MbsTyEOT
jvEi2YPy8SZganNE4rVemIObqUxbuOy3KJ7wg6Mamm1NPBFWHdsnpxg/XHecHBEz
cEcPuKN/gvQwCiYWALiML/+PRje9tPZph4cvtCjzdqLeDNYtE3fCAbe5o60hZBzt
se+eWib89P9p1RjZd9KEcLrNRgt91Aw/ueJN0Id+kvUnHa74WVf9mussl9+K8Syw
Xydl/DzSrmeC2SdxX2sXUmUR009zZvHlArr/cfOJWq6ryBb6dd289fMo03DWJODx
QB9JD/gNzd7n5rsj+vbQRs/bQa0MykNAwpQDHMopqavWEz0Ax603keUZip+UxDpN
eUHaRasXxRmBOTsSpgZvsstQV91cn7xMXYRJZhaito2XwZJUG8IV7W2dnx87LfWR
p+iolZE5U5J07KuWbhnbFwXRZtIv0twAQgu1jeHBOD2tzsppi4czxbsZcbwgA3n4
27Y6bG9aGMTI6r3fk837ufJoOHX6aEiuMcpqy1MU8trF4dWWaxuoT6EOFJ+GSPK/
cQ2fofzoCVYykab+CLRyUwSQAxjuVDQS3yc6AaeZJt/jY+7/NHPyj6wjiYc3XchP
F6mX3R1WMLEeox45LyeudPTqfokGzzqpP2Rb++YjtjlTdJTlXBUdWxH4zDFuzQBU
sfBacw3h2JXKRfPrytM/gbLLg/HM9lCfnwqwbvvU0GrhVhtqJoCpFA+ILys5Fxvw
LWKNGHsJXWHUD1ZzVN79+GCvkzZCEu12dvFxhePzqUEyHnkEmx8VJuaLNhEOk6ca
W2cr6wMXw0CjNznnNr7x31rEnmoXYOO1fa0AMYTlA5SIcY2CW9Ia/RDOOYQsQ4Nq
EHacRBTNI3pEFZbTy/HNEq7pMIGvo7IdmtKyi6JD1UWT2brCw40PVEvf4YhoncnM
FpLwN+uuAzv88lmLPvizKKUBv/v8KyNmO8Pz+PwG0P42ZDXdLgceBW6peODAPNEO
hxeXXascXZB9jfgQIVF+oAZvpYCTrlsaCWSE4S3EGR7YbySJBY8hYDoRsQG4RMwb
g9ZPqW8YY4vmFxcQWTbm5S/6wyN0KXN0dKxP7xjQHs995jeujIBb0Uq4IiDWK22q
1SVp406WUjonnydIGpFQX/gtmQ+WzJPtlfu7jB+lyCpEEZBQ8A3YfXH8swRx11Vc
kx6hl74qMrvgLTzoH7TVlnzD+MXo7E4ciwwa4V97HRQ1ArykzaNexIbhE/+KmvUj
uUYbwLQgj0evUKMw4j71KYKRrv5ruDFq02LQha6o9Gemm9sSWQrJvWPrQCfHXVJX
CsHHBM4FqdDPOuuazyFWhSwgrvX8ixWKfwU1wNNqx1xVmvpurC+OF8KNaUxrpZ7/
5cjvTtv842NAjFskpHQ/WuCKHB2mgLnPBoUvk61RSnihol073LZolXYmD2TjEdb1
6rtnpWaYWXnCuzWdW/i9v27DWSX6VQBDcdkD8GPKyeGuzNlcmuyTmk3+LSKjKlbf
h2cX0k2bArb/419OrD3/ABeEmVIf+S+C1ZULy+kjzn3suCkVCGRqebX1J6OorSkm
cQ4/YBf5sknxixKCkoGe7hyvUnEn82958sndwF6HgNQpFBqTisY5gtpePpjo8BPj
WovOGjHDZgtyH64FGLGWo1LXPYHDh4G7ZkEnEIfXm3kmw8EiX2rFVDI8U0xJ8ASV
YYjqAHBrwCVnMhn8aMFizpKjL5b70+/ODPJgzw08BenbWhUQt0dH7cSqIbCnyWBX
F6B7fTt8qRkuQuH5pyGde0RAZqjSGgdxuUByD5Q1FyhepJkictBZy3b4THQ7cRxj
L6m41h3G/2xM2g2jMbm12CfowRpLcQzqwns25JgYDY7Ni0AiauyceKj5FVc4B2lB
hcgbJRdu5SRPMmScazCU3UecNtQDY7lXHN12CcPUypVHd52TF5SMAB5VK4ypJ1w/
r1eQ0joG9MfXX9kMdaeJ3uudK6GcXszgh7Sf1CcwbjAxDW1AMSeYA7nUC2W8tini
o/KPDCdIwoHsSGirEELa0H76Y244cBKSzlB1pgA9kYN2gF06XWFNnwEC1mACaR6E
Q4w7VNmsahI0IkoAEi630IImxfbLZQEw+OAyJhKxiPDNnkVneJDo2+TnTvOR8VV1
s+NrOY9MInNwJ/QlZ2V41JEDzvzzns8jJaU9xj4cGP04ZD2qAS9AZ20ofy/6UBAu
ithc/o8I4fMjBJ8wX3oHXsQr4T4JnwFZmFoGxzRxqEuuILY6VcfnsHlzlZNw/ftq
hSmfLWqvOpLlTXXwi4Is94X78EFmg/vlC4tHt99Le0gTtmQEf3KkSPYgWRYRstzI
TS3XrttNkb1iOYFaSPF7VFxtH/TzLtks9HIlrsF4l9qmh+OuT8JsCKhqp55kfdk3
oSQ0nt244+sDq2UljLJB7Q7RYjTL4p+A1valtG7FLC0m0eRqbNE6ILxMgTyGgzx7
/+68zVRDXpBEhXHDGw2wp5bvPjUGwkWFJn1QdBueK15EF3LuIRqkzzrVyk4o8Vt0
9lY+0oIR9cyqc/nOJbzqRu/4PvOushMiVxjqD0k8G11HyIMN6zjFl0rvmJDKedR6
zuZ21QxyAXC01j4s3/Ghg7/md6zQDfQzrKs7svpHTgkACENUV0WZoTZcIV8bmFDR
hJDiMu09itRHYuQ/UE366tKjZVASoVJ7Ze2XmOO2QDimbRo8tNviS8BKueS7G1Qk
mVYMoobm+ghTgTByPJAuAXlIAn4CQVRvIWTdbd6U5lvjuDOKN8UQC41UkERvFras
F4GYJERXSDhi2rDunjz97c4yLSMHdE5+La1SxpF1h1gG+Eabmmm/8dqQimAQqJ5/
y8ZUo2ln5fqG/qmS2IDde4zXikL4rDpt1C4E4iVIKJ9PxbOd2HtQitcwbWZJwFjz
Ub+Yiu0RRosoxLYWPxUGdzBJxNVSVj1aeXhDdl9g7s7jBqJyge6nsgL4gDJz0aRp
lKCcmleBey0lDMqVkTAoE8NAmECeWlBuPPB0HZ2ukd3oycd+/tws4ohcG+XiF9zc
mOKS1/y9jkHNE90okuFvbDi+k7Ab5BhPzGTBTUa8ZVBpZHNC7htMylca6kFkndC8
H6vQw6Wo7GP3j/h+0XLpnrQoieeBfV8tOWs761g8jHanSmgLJ6VhARn3QAUTK5m6
3oKOfbagk5Fc1PfEPVeS+88030xJbzHMnZbk0CeVJn7IqHzNGY+O/BQB4UIyYLW2
OYttuzjiQ8oUVOltYPiLKTXeQETrPL7JffcHOcj4kJq/54+JlhM0wtLo8eLEfUMw
X2UfesSDIchc3T7b84ZU9hdYUdH1zFyUSxG7c2OCTBOZvyeLZYiG4uYVamNg7izN
jGFEiqVAFRAiDK0jiCQIqC0WGD+ikcKgGFnPGlMO/A70cFwoftiAE6L/QYopxscG
zI61f6dVD+2XjMfm7tWKoXt1zmV9mRYUFLvJTswwX1nuWE8pgiURVrKQ8WolBzp4
M6eEEw/MDzD5TRcnsAYiptJdtvKmvMXWgMIqWMxK9Hi+ZkFqLr7u0cSrVinR6AFk
TJjk5pq7ctHveEvefA4BrhdEKJ2SdKEeE87hqJ+ejR4syonwGxm0pRS8rKXv7G+0
C3mxuK3LrTrTQK1Pev3ykfAwuEO46WErkoVxcfZZxhVnSFoPPRb8cxXEVhdO4C4z
eJwJsjwQqEgLWLbhfG22zGNRTo7E/PtojAuTM2mkXht6S+9xWDQXK7SDn7QontgI
2iSblzfP2NsPLICfZ5psIJ0O8lV0q4Ju3g3gO0KFbVM3NdmHHhAz9vR0RJVINwYu
IXWiStcvy9SdfGTxNYUHoKSoCtS8Eyp+qlIDgz6oS3KSaW/1QPmhNR+ogsbtc9oI
LWOrOP2HL+xwNjb5ePf7ZNOylMEuTKyX+kpD9iS/ncE1X+rsn/NV/PZfKcjSD244
1Wqu6/BW84dHJ7a4sngvGMu4S19cE8ZzjJMPt5bZz9XicJmnDzPdAoRWkNadOsRf
kJMKzI4MRBsPBBpRWCBoxkEkTJhhXbnFsH9DJAlp9QK4aNZqfwpJIgJHi56UFb+q
g4zlrzho4YoovEeY4eIRd9MixwOpQSeYWyy6e7P8EZaUEIZl6/Bjfif3Z/tzQZab
ZUyVzdSRWExtGt5ePgHclnj1tr4/mLIhizHmmDjn5+2i6NM6COSZuami0P+3TLf2
9hojefi5UbHyyJGRaqhe+Md9S0/me15UDi3rWmJnOg5bCxht7SKaWatW6/I9bkn6
uBizcEJVs0qF1oGxydEdbrY+R2HFPVdxXNGZocFaz7Si5JaALO4IJhMhMGwyjwCw
BR0U5i/+ADXFbcAJr5Utw/nPpUoVZ9xeJfjeOggk9xifDX/4uOyIK2dpl16/20sq
DCEoeuWLJZ8ubINoGEId36oQjx1eQwFhIquu163uQdIRtqi6GyxvSRqtJBAoTGWw
YZ7dep8fYwclQGyVUexEnnQbsfx5ZQcwXJ+e+dokYYtCjkviEInmteKNJHRYFjAB
kVzHUL7I4arJskYxM0B7IqKiKzcmFVdRH8FNSzNv2fjV5szrjRJK7V6lAEb9UyCK
hlZDyFkFBl4Mgjcl86zoJl0XPXibbyWGKsYqjxiNfCbysBIby2NDfRneEGmDNJ5e
CAsW6qar1QOf5OIEtrNxVIH57Njd6eZ7fAyyzx7brpDcz7DGhLrisU6+fwMIsG9p
ZZwp7xFtyTfyjTQUQQIxKuKTd37Ks7ua+DKXh7K6LySWXQcNqP6U9QCQ0iJNebn2
EhFr3lbul9sCiqW5vWpOmeICmFoO2vt/QoY/DnVQscLcrLQxYwaxsT41p6mDdX5J
YkAB6/tOVK82VuYeLO7hSYUDDnJXml0tBPA0eMdkVB7gDR6t8a+ndsxS4dnEvOZj
jy+dPemgkOcHmgNvZYrnlMP/YFSqJFcZP/bHSQ5d/SoLRU1/qBJJZqYrDZnyPPtT
jFAM1zaOaHjuaVC7Im4r9004cS0vep46G7oW8sQZpgyN0jaPOGJGGxY9TMAt/p/f
/Q1wCq8RGxuDTr6J2gOWwXl0m5DtPDhchtw0We+0nBZf8Apxk3DQ5lXek//48Gzy
vp/uHfNJQM8BS/UUtjZFwwwMAAB8JbDDO/9n0EmPkkrXtUNTSL1ERvjpgqs3dIop
/RWwRwSd164Cp++87nBpSV7JaV18+6pEFlmrb3c9DhelwUofNuply/L3q4XvMRtX
MjpvYtZp+OBBHwvMY7KeeTfS4AVPqWuw32T930jgfUd9C2BURfoZB87cKmoTBhR/
xZQRVmwJ08qIIBvDCgl5w09HiMLIdQWhEg5g0eK/arE3/4zC2JcUMgqsxVrFggVK
uy4Re8+1xKf/5XeJU8ns0nQovJYW3timNdIs3HiWPUD4tGP+mJUl0vkdOYPw57J5
V3Ufoop9IRlXcskmNHv86MIxuFyqPAL+JqE/eMCRygTSpBNx+Er/AmhH9gdOm2II
ICA+IjtC3CrdCux+puQmhe9d0hjlBI8IpUxAn0smTa0GRC+MI7CwNNPGTmhJCWy0
Nrn+Xl7UcKCkD7x+dnCWWQfgR1VPz0ggBDq74DmviXYR2CbBupqzYf+xMhWNT4aF
wx6ZPr0WizVEIZTu2VwSG4iz8T/Jf/6CvQpC/Cb9/RjEc7l2UXC8sYLjc1DZMI3z
c57xI333Q9aOrbP9JO+iJdAkzdXeEdKnl6wfHogd08UUGIttVuiXjcpl6os8M3Mm
Rdctd97gv1IGugcMzwGq9eUQa87vpLHM04XbxXwqjiAVkBKosnH0wEDJ+kHbt5By
kJL3ZhXIQ2G4SWD4b4w/YMwPQInUhQ8yPCcZpdbvpY/vU0ShPyYMf7E5+t1vFnBA
Qtu+jHPLmliWSQNdMbP+F4fCZixwjb5mevMozAwTIHS89sEkvcQL8L47Ac5apZum
MeJnHS3/pGMKUpxCfllBrF/URlB1MouIrkFu/SUnJzGR+7bqHeMjGShMwCKtW6ox
1+BX+FK4/XF5zKbyeyzdR2BACPNZ00f1bRcKcJc1DXxTamy6QZLdfJyC5KDCTNay
RWymCEkj66UxVfWrdT7CYo5le7RqN7NnzlJNiMTxyNPs0113UKm1dBbe+hURfI5a
2Nj3O4TNarIvlXSyE9WWjeFa0kYdtfsiyGc824jH63ULfhjszpnpVCFd4ZtbM6kq
M6JpJVzfLy3gRGyePeI81RQrQILsKGPyt2IRX7AAhoNL5eu8EFy3Mnkk21H0t/7m
fRnMNNlYdCYGHvIo8p8OFRMgfYVeIR7tPWa15I13FXIMqA+JzirEIxKDJDf3fIJq
G18RSyCVdm/ARreCkkF9ZnVD5zOftoWNHGYUWVPqbR3f8fS6de4UyzBnbP4ol9oL
JrOXCYkhKi8Z07MZran/BdDaXadROJfJpOWuWzI9ecA8DDKa3X/NLRsDFeY07Rqv
oE64++Wus8gyBi/H9RuIEWEX0T+fdgbA3P4++xjhlCIwZbA8tW/x/127MXiYy2x6
IabkrIpK7Pzz1Xl1SgaUlcdNdD9ahHKYjGZ1wRKcA+38AMX0nHT47oHuNcAa1yo8
ajHOD70mto07Ik8hSuNejrjYFyy/6o81p8nHgQh0tcZIV3vFiYhzj7iBioCwzEup
n4rM/H3ard3kq7mzm8Hz+URFjoW0+gteal2NtYTgGg0YHJ1Z5QtEq/aWWtiMq0Mk
9vYKPAhpFwvyb+lJ704+hraZIrAwTbeZoKqxHeUjDMhHO1zQr0vshLdGh4hJOCPI
13RX67q/wPaFnTEbB+ZluXlrIXjWt1F4cx0FJwOCY3IJLJb03fIPBEbhn40Fv2q9
6/ago0nVhAXQFlwbBUntbd/9B2H4XM936dRJuyKV62LYLv/LarycjzBWmtTASvaL
gHLijwhNDGEJqJ3vCFmMBDkpaGyLOseZIgvArpwded/AEG1kD7Bnm2kC88tJNVn4
//gz4NUhN+RpkeMXPYc6XMSFXNun5LvLj2nyZVpWNznHgdt+kTsd2hVbnsXcwDV7
0NHoNQP8wo5omocGrnuNU6Gu7SvflGhcCB7fCtzN2tgooz+xDn971wp/HQOGUhrD
/Q2J9wNz+ofE9mgvBYwD3vdZWaEEb367jZo2uk1bCoTYaaPnhm//JK8CnMYi4VZw
ueq5CKyfxcurLixZNG9YVCNDuDBeeo6WigqVsypjl+InSFNsDFnb6/asMKjvG/bj
l79yqfFriE97PVkKqhO6JTS2T43VGcYAhjy8gfnXet3VVyUQnKHC7Bq1ZR4eiw7o
C1O//hYc0o6xO1IG7tji8xPT8+qRIVmvgxfEgLmZNXAJkR9sUoEqFXGGoy+200sb
LYdCEA7XUciZnPwsuxALExIhjDcrECJ4aYQX7BAUubzPodEpTYVl1b9zH2QrTBIc
fkSRWzupJEvqFOoF4Q09tw0SOxpfWdaOt088BTZBm8apvayCfz0PUtzCR0K3rdPe
pqKJTNzn7YmYtZQumq7bkhyW6NrWZo/QtaA6LKWYLtRJq3S3sFmaEeKr82yLa0tN
p6qqvJntMW5wKCqMyvOHv7nDHnbWIR0Fh6uqVsyQHeKZEHYGi1QTDg17+rIiC6rr
mIJ2d3rOgIZ+z332/pgXrSIHXgP7/cbApVDLPdxyjQkBW7m7D68NLDt7nGs9u4yy
CkXLbo/Mfx9YuAnTxLa548tJm+K2BN93rethKQ3E/6AJ+eoelpe/eJPRYllRqs97
m4tvU/ECkd1iOGTKc8VB13sGgHNsCq4Ls5TUo0+R2kNzoSY3DInpmvqmwlnokred
yobZzIOFSea6rlh+FRHPN2euMR3V0nThgCfEzvux8A94VgzgUbUXGRhovPDg+b2i
ENpxsjAQ48SembmbGAI6ZAIsr51Bfu5BkaudmT82LhKOBI3ebQBqx0Z/UnRpDvY6
BYFNYli8ORI43+RlqbCIrEviWgnWnLMukiBOSwDyiQe0p9NwMYEUja4he5u83oHn
UiNr+RN6zTxOsXiHcCaZThVDnlIGl3jpP5I//u9Cae+panQ2JsU4c0liTU5kk3sd
9hMGAjxmaCX19MJ2PMoInlAFaWte+9MVeUGRhkKASBf7WRjInFyhKD//tbpWPNVz
jW6BeOJ1JWhLybV4CQodCIt7ZgP1Zx7Ej9L5We/UgFdqa4bB8yCqHmSMay1o4jbA
YCYhBRLRwJRyYR//LM/TzQ2VhIY+Q9S1uctzXGcja/CvKP+uV/zvydsW9TAchNFD
Ul9buh4lVRcHlPQABNw7gloljCJG0olg4F4iQhuQiuibHlmgRPhbEeLu5PiN4BKH
Wwn36ep0ShByH9QzJy69n0RJz7VHo5bitOfnxS3h91vC5QLmy6VMHAjhSQqB48G/
6Aac+QXGbLZKqngHaUyXh+UZgDFyVFXlwqsiCKBJx93T50Q4ib0yyUmsl7nJ0y5J
JDJBXOYCZWI01ZQQs6rrDuALGhZQ3zYjJshJCh/O2Gq4rXESY/6EdWJvgMttDyJm
CRKzQLaDLoGB6/VigWa/a8JSeCKsz5bK61v4y+E+0oQfrOiK9+mhlH2xnG+YKuiA
BDjMIXxyzWFF0RtFlrgq0R8G8BF+OByuY9gLq7w36ZK6QMs2dC5KU0omLYdVfYJO
8lyuwMv6+nu6Pdmh8kVy13MURpqtmvw9RB+efxutCISZvVfFH43xhcKNZbPnM5qk
aWcMknsFagToqb/BXfTtlSxqern3/I5Q19AjIXk8U2VA2v/SLvsNDRSVABn4yAY5
pZOam/xhzd5fRYo+6PaMUI4TqZd0rT8RpUOlMm8Pm1E2H5rRc3QOvyvV/Ci4iJJE
/yap5koTmqpafk92BUCYY52VUUaurEzwD5ydJD/LC4VDegjoqXsZmQv1uHWPjnx8
QweMxtru01pANM8D/51lf4PQotlZR4aUWiw07nERYo3GlLhmDyTUgTMwj9sQVI2z
IiRueM+h+B/FjxeDFCbBfG9gB0E+Taie3Gg4z/lUVt/W1edLn3iOk3Cn00iTRvrh
DlwszYmNYt+qjN2ILyzGEmij9zmPZzSImdb1PuXYh/DjuvNX0iR89g03phKfl3+W
YLzrppNl4BXvL1qGvy2QNNuB7jDkrJjxFll76tokenglSoJ0FMJ5es+l1ajKaXyo
WKdZ2kuxf+OKqquuorPAAwd4Rm82gjgH92rJqO7DziTt0REUbnjbhQLgyOMjkOs6
NN/Hn6Ym+egdPI9OUoHhGkikSWc8dKeGocXum7ZM8Xe6cWFq2Mss7P14kpRIyyd8
Z7xR6Kqs+/REikRQeY/GTfRx1jS6V1hItKnh1ExNgpjqHtLdXAaN3KBlcVhzdvez
WnA4S5BCorjjPGwvW0wFLWFrzIMz/1Q0s7UAm3e4pFIg0u8fIqIgVM0rkrHa6hZF
USMQPhnwiW2Dbrnr1ovrey+8+FpUUQa8YoMheJkLE3+E0cIddYtEtYcrUwTocp63
/FAZZQXCDBGYwrUf28xIBRu7elvtFfjXFc6M0PMGa9iQ/OeUTTtujs8SY/vkXYqG
1Pp2oKLHDAOjhmRNpKmb8WB0AjPxNiOor9d2McSAwhhDAwm31lwkQep7mt91/j+J
JrfLRxWybRGltd/Cp3/4y0oHwu3bQBtiXFVfjrsUXj/5vLnLczmLBWDX1zhkDzdr
6Yx9X8ZHN3I/Zm+jqHxsWn3mys5M2AExStCe3Ew+e2sPcJorAVPtDG4ATRWML8h8
Rh1Cw58HuaXIKGQSPDDDA2ZjUyR7+Nv+vwBz5gPAvoIJ67MCkou+ptmtUQwv+cr/
qM/3ENmEgBc10kWeZbNgGT75zfMyork3CrlDNPygyZ5Dk25PFxGn3nbHupvd7OCa
Z/REGWjitIxWNsMmIS1didQ6wxh5pbGGule6MWexXfWugqzv4CPIIFcnPtyEdpHp
b61ahb5T6s7+yTnjph68rndLZcp60XRX6KIeFbtleRj7AjJ2xk7MaEAXiXMsB8SW
y3oFiOPCyjWYEpoBc9Hswxsuk2X4ZBjG34N/7NFwyb4Nb8wbUDjpZs5NF3ygB7NI
2qJ1bPdX+qYYijc+ZidMwn6Ydac/lPqBKSazWFLpnZJzg4TEJA1b7nkcXrSfILuZ
KfGvK+IMxIz5ko6mXHr3WhCS1GlvwVVxyhAwKxsh0D7te0oIzxnCqjNPvnluw5MW
+QiISmZmlGjwSi3Wrk5EhLajpTdUg4ecqlYLrDM7rayQlFQbHzuERSuXCpCUwvkH
nMJ73qBjYbMLqnTrFAg82YEnrsKbMLGtyzqCW1kKQyhUX6wl7/BTNbfRGlH5+UT7
iau14wMBkHRoR8c0jdal2oSdP88wiN9v7UcmXmT8fHQEzxpJVEkB0bf0I3AI3X2z
2dCRhP8C4jtTV1E5UQU7mJyqcLN8xDj/dFDly5XW4zzTOpzcpM3c1GXMhVh5Xf4K
+RiOvLCo4rgyy1qd78DHwoeiuL1XPNmZxFEs+XWtVE/CMMxYlOKqwITSKPlL0JGD
OxrcvHrgrMEEslM4xNrPaPi6HLrogXizv8Mk32d4XWogQoPFuAAOalxeiNiwxW+J
SrJ1IhsxdMPZtaZNxHFyTdLxCVTCq6OjME+LlSBnJPLcBckcyrSgBKz3jQ4G22Ii
ajXASuaA/CJZaNs4y3gsM5YDqw7B9z4uwZXMsUlsTdqO2fyN5NWKawI0HtHeMF1N
ci0ImqerladtYXSskFyqgw+otTF/yq6+ht7tGFaclpdOknS9cmO0frshJB6gkT+l
9fAVh0k9gKTI0NWF9b3GHL3NzrrrltdWGmPJpqj1aIgraiFCtmxGyexNIFfdmpMx
rfNHLyI3if9oxaLnN45O14LHATXLdXZb2twGqOOwtWAuGmCBt/2I1BKaLT8gd7xH
h3DMx0aMBpSQLRJeFkhFLEUCGRrkp1R9RrYe0lEKdyKCg7cq9oII8MejZYSHXAw4
X92VSNXRAPT+OR3C/GzgYFOQeKV02trAkkj+bfy4ZQ2ryS2/1CwcKFlz1K157tdz
3eyTU2K0sDKrfDkiP0wVc/AlOafcmxw+MdBQM8PBss1yoJOp7cEG2mJj2rkeJeSs
6NCg+7f8dKYPx7Pyo6ypZjgYz6Gf+7mZgxR8Iva3r6jRHiFkZHurusFEYzgSvenJ
uzHUSMiS2rQdel/wZQogzSF9+F7zFiP8t9sUy0j1jE0juqd/WiNOzZuxfXnpknZA
pc+W2KnaIvodDx97ZctUrOa+ZIv+e8BOBIxSABZKzYokZ2kKWh9lJVQFFd33qynv
7LnGPM9FAfYtK/BtycxOlgXuHv4DKyMhZhdUv6fGCWkovQxlARV0QEi8dJdRUVEB
eHQ02XzHyZD/xLiLc9vzANseDOzmB/ECpGd7KxnMrjH+xbsq6A3Kbe0p10G9nHf3
j+zh8M7d3DrmYZti6iMqOEmJB/Mzeq+DvGM1wzQ8we46+N3CQOTyL6qdq9vOMfpu
dkVQEy6AaYHXxORvnTQGeLatkQqwJ+6fuSmEGCnuUjc7TWh9QYaB+gr9JjB+Q2AZ
E69TOYYZjj8Z2Q2TVEAm5v9kY3hdOdHS//ZtTDUBdk4wjxHHwx86xv330tRwtgvU
Z7ZaSJjQ1wM96JqCHsX+Ar9i79z4PeU2tgYPKFW7MXZSAnZWsS3y2yHZQsy3brhG
ROub7XYCGtqSQBQTHWqrEzOorHgow2AlErGzuF/Nl0IimbGj1Y848bzLdn/KwIIr
uDiK1pvyCeNloJHao0e09LTCRCxxKO5l/h4p8aNou6yP46zmUDI8Nq6T+V16nRa4
sDLYi9oM3tsPojlJJ303tb3Kuc+w5uybK6llxrjOoIZ3PA8+ieKypZ34pX1IPUXr
CFcWjzqgFsKLJubVBaso+EHJzl2PJKuKDRXEGX14FU0e9vbszFQhuArWWy8cZIvM
65+955fUVHvt6HfNF5E25S8FqkL4WU+VkEDZ7pP+FA9rzoZQnxKhQ3BaUKP7DX06
v8EKn4wd6Bnqbym19UNAe+J9vyoTiIUb57Z8hVP0B6XB8J75/9qzUTP/lT4MI2rr
W3qK4V/BtWoFAeo0YKH+phieFKYjX2ZForAbMKUKyio/mKnEGUNTuMcvETCyZ/ve
fM9Zr2UvauZYdE7qPGlN5IkHx0sxHStNVipLshZn+cy+TphVG4l6Y7ddWFQFhJEF
a6AeObGeAbLKSoo1tkaXbDRa/QvpD0RywjEEfJAEP3J0TOd9agQ/zUO6yj9A0XhL
qMJIEdcx8gc1pzS1hm5rxtOceBUzfnrCkKYlhaK7cgbkkuw633emhffN/9qy0NaO
YlDs+0RPDngKn3sfa83oF9EAkMYs4kItjrBeTxrgUJ3XFdbGNeg6bXhAND98wRdh
IkVp+r6Kuz+JK2uakHJqFSSPUH4nrgO3DlBIEo3toelxQddkDo1BT3JMxdD0PFtJ
pkT0Zk8ukNd/vEvIygfEIhfYxKoO4LJKh1HnwnDCjtc5D+yNpmJdqslGM0Q1+xT4
RyjOPavkx4J3x3SzhsQRzJla4kFEn/NuvV6ljSX1NMC4JuXqibNfSMTN+VHBimcB
QCQ041fZe2L5XAvv6hD/QeZ3hOnIOUpvUBEtdR0UffRS0HJutZEg/wW1XJrY1Zhd
kbBjvRBFFzb3NffZVAdhFrbx5kOuj2GHEkJz2C4ZJMp27dBhLAyhqB7XsVgn6fPb
bIQyIzZFjpd9GdO4jA7Fj+wP2/QKOIjXjw02qqjgnGlVM4FJtQFcHliJO+z+D8zj
BbGjkdQ5XJbwqdXcFwzQOOU5VjNzCJPVeXvwAwY6Ehnx0cQoaxuy3rx5fUl4Lnx3
0QBwiq6FBex4c8Bo2f2nQW8/kFrvGCswgIM8bQwqC6Kc6d/VUu1PEhc8ltZFfghh
rNlsTp1Le2NzBCkFOx15Xfu7xYqXHQP1UFf8jaV6ZXpmtqeY8LpWa00+WBWRi+4n
CK79TiLvJlLiAGyAnSPiNh9zZLXtM4FxuJKgD9/OAw+hFpvG0okBPLhSs/N2aon6
bkYGu0IZ/23KsNtAesCMSlZcdFCsGN4EklQJ9OlIghpZD+Z0UggGv2aVr/CW9nOo
Hs4Vnj+wr2JSxQytZHMUO0UJhtvrDCctJhsM0j0ofT3tsdL0vbhqtF7i+YE7Nd2k
zALIUdT7tzZQRkJMHPyYfBHJoYKUQksKuGBW2T8PyxgD5gxEfM0QvTTvfzm02Rmw
FySYtyixMvpGmgAv6EpzS2HuKKLJcPY7Fh3fb/MRL6dxAd0Q1PvWfgjr/ouWzdpy
ReV1OzVfH1tDTVxt7+yhSBft2uBI8S9giMrtDFAp7deBILVzPyM6nJw++g7d+lkg
JKyFrO262MAoZa32UtI+vQK6guBDs1YWbglEhcT60ZRqozxBdQnXSOWtN8mS+7TQ
MVoynDNcFxTU0RKy0nMkhGDtrDlHB7bI8rbjRSmhszKWdoQ+sVEamES7NoEeS9zu
ZglllBQDa97abjpuOaw0lnr+dJ09bwRdallZvyqiW0IE0OR6EWsSEFRB8mLFUwyZ
2I6IYYSRmri6p+G6fX7zzCC7QnNMGDgg8RQRvEVi2QtGQXQEIAWvk8vHZ5VLQORk
gVLhybPrAK/kUT5yU6NIJahTyT+v8K4kS0ZHDslZAxsJOZjA6E/FVTo0FG2V9I61
Pkl/DWTvC34u1yNa6HnKW7afiU1lN08D7CExWjOlJUOanyxGsEqKigfs64C3xmCs
CvGKexitv1fR5O8BQ663hpRkM7K6/pZIInBK/t6NN4XIUAhD9syjA0ADCIEqPUhb
VnHwFnEmmV67lvfQ42StYngdCrofKmC+WjfBm9Zkq61Bfd/z3mbhVAL6x/TgvIMY
IP967XsBEuue5VcmKGB3DkYVO16kb31IULyiPlGXtuZL+rsjZZ9Y9ALPXSqd7tlr
/iS9rXhc4GPIMVbwGtnFmJejL9sn8Z1tzy2cgcXdE7iSCYElIB7EXFqM7zPeFxgR
pRqnhKXiU89Pz4IliVK37atYKmn85fRWs6Gj6dFOo6NLS68h2UVSMkam1+r4TAqd
bwgqDGJyMzcmRwePl4li/JWmOc0+WMU9uZeh/HA93gKQ+kPJbWuAnIQMsjQkWYqw
Fg9D69n/E3k6B+t6QIUgnqmFRmiPkuHaUY1taMgfrPV6w8S3CNwZpI1h8UgOIWcE
ZCiERkXVcsmWYGEmYGVIU4jIxVpZmBpTr8iyN4HNOMZ+B38wg1uVDxYQrtmyLluL
PBzuuop/LxZFF3k7D6zwGs14/awm/MifKaihSm9NXtUGI5nLjT6MeMv9QAf0ZWwb
DT48+UdPvGU4gRRIacFZ9WtrzwRUZlWSfoxJw6JRaAN1w7BQbJjWH9RNMctnKR8W
2KLAwlmTGqwwXJfR3wPKWCyErRPolPttLQjOIRMhfFVEFGRxQBacoKw4ca/2eDh7
SE0roY6HlkmQjcVHPgpR667+D4/37BkM+f+L+wbp8+klcwXObtdhWIk1q+YWMqeY
72tD350FN82wMaSSEwhm/MblMu7x6YONM1XIISXMSI0aKkLgVuXCEGTb/laYZXcr
mNj5joYvXCI9dm6StRC1iSilrR+2rBe6W4BUBDjEWbkN9K9H3UN3yI4Qk9Niv2E5
1a6dWXXVNN0CbpCMM5Sa7vqNEqznYS5PW/dqAw5pzlAv1KkEKCafIhUHU9L1dxX8
cheF92Q8NVhMaWaX2A/lxOTa+HZwM1SOQUlKScpu8s9RtRS5CRoIMpxZBEjct62N
QA1eD4xdl0+Wu8ZctjhnluBgnmc1HJuaUqQAWYo+btdLL512j+m4y3mXKGKKUerv
U5J3WFjEI++E5Ga7jCh/I2ZSHd2D9kkuLyzi25hXDax/+jdAUF/QUW5HSmzEMdC9
KC7NaJyzC/VHGj/YyiiQcdBQ2sRJEMEvbZfRR7Acw6EIEriHJ0EQzEThklveAxK4
JWJSVNX8Lw9j69Zos5WleF4ZCXd1NYc/OJh9v2p1CK9Koti0h0AABJxY6DoV/2OA
7/ou8x9EXLlOHC5XoiZM2NLNzEa3jw95ZPfsbS7MndoGd3qWm711qsZIcuUP0ZT+
r3IPo9nFtunjwaElkDJch7WCX6nEDBvVBlKmccf82znVDG4J8pR7Y+koictECluY
Ynw3H9Ai3+qyVA7LApe9ShcVmkrGRNNwZ2yCQILIPm01aGnnoPa2dt64nzEUU1yF
tnmn65yinNSeZu/qkK5TejDc8+zYAP1o+3N1nomnBKCepmZCInT/V5caPTVtI5Vb
+9uHPvgHGWsfTF9Zn+xEUYOuK8u1QpoRHdj7IcQUwemCWxgXXOSxNCkHYvKccq0c
VRS7HiyEMkZT6O3wWuzcgAqn0fyFRMwfwnplAmBsYB/YPfQFP3xw81jnu40JV9G+
RQfiLuM9cvv0nokKIzRyAJuGyNWNvOwZKckgG5E1+epvGTSo+/Ip9QcmKbDmbYT+
TrC/GDNEko9vI8uB3SfAtCZldRb7mN15KduEDoeYeRfXgBMAWcCy7nhTRVzZdnHo
CI4i4ALidXjBsQSKj/7jhIJPey014XJgjsK6YsLmXMPIS0c3KN9TvEYRyNdhDQPH
BeE8+w0zKIEpofNxA+2xSxGN3zvN8X3DXW4OP3FvIf43QX0BGeP5uqZrCkgKG4bH
4j8hPlC7bHYHE29G3BKw1ZshS3zr3AubjojHjoQM5DaM+IMPCImVlJ84sFRutV5H
H5jjAjf1FuuFA3qEzgb24zXCcKlc+5gkANbYusRs6RFq+lD3MpOldjW+8EnsC35d
ksNHwWyvNiYcWMrB0KS8u0+eE78MlvYQa9VROmYAIydiS72dHgFR88YxAwGXu9UX
Ntfi1daL8oyAaOWRlTRzZ8qgPMwhAl7pXe08f80U2uSn8zDOPNxdwQA0sfN5Xd13
WRKvvSRLJ1sc0ZdXtKOWjhJD36JVgip59oyCJJmsCwF9g4SFQ0PIYrIVZfwX1UoL
hUpFRnZgtDmb4HFjDYkrrKTNjNNB2kpapltVFb+EVI7rspXPZd9Hu9uTPSgqmw/P
i9Y80QQPL+ta0m2DDZpUxq+oVfNRoWwM+DYVLBBclb0TLjJjsLrtBZdMXv9yXqKx
3z9KPl6v4GuJtXwOlvyjxn4uetBc7qWpeq3icqrQ/GgzCXb8gbskYQbcEVj27DXt
CtiJs2zEafdrHlTs104R0FmHHzh+4sMWYyQMl8bB8yFzO/XtFDXPKRfhx/N0wsq+
PMA/dId3MqrFepmPM7L5BLbU8OxIAKUgSd/PBJ6carAO8c50D1XkcicKPttVk5GQ
Jl/8PF31y2DJ33N/n2Hl6XPZ3lTpNa0ZU15L9pNfLlduFGlhpI/154vDz1sSb3y0
B3I70xmV/6fRzDLPl0K/+q8o9xkKzcY8JSQSLVIAS2WbbK99c4B6bJatcdMfhGq3
XEqPWAJNdMzLTntsrxVvi65f1mkFhWKo1/Ni9tXSsK03CFVQmccS0obemhPdQGhs
JKhjtkWHvUrnhdaR/RMVhKQn3jzhTJmkwVfom2Xo2YI3RafjWJHr6V50KSXTKX51
6ytsICXw+fvY3LsiBrIKgVvoxCG6jezApTLXTi4JWHQY45WB/cDeQTE59lCixB/l
iRWm8DeQN898sWF4E902vjmQyqKvc9ESZsWOcYGyRxIE+ElF3giDz6PgMIEaMU6a
6LxQN9QcfzR8J2PAVj9VUbAeoYAhXc6ziGe20dIQ9Je1ied1ai3JusZ5oYSV88Hd
PWaq3Js8xr/5g1GWOmKBkJLQErl8E9MtWO2ntrpk99/YvScAlvdubY8g1yr4yv2B
tewFRoLAch8gq7hzoNj91FQovh12RykKXRiDfoRwKX6KBjjsA5FpGr9QQFmEddb9
P+T0wu4KrXxERzbmadAG6dqZ5D01QB1LFNehD5W2k2OPiEKz3HSQCYVGNt2IEQ+s
rLZrHAReTW8H0BH6XE2e0wAf1Kf78FVoTngti7BnnH6DuNR2FnFIpNnuCmj467i0
4Ciuww4JVPvvvjFXE+rbfABLi/8c0qmObnnXcjSCSRdj/XdzHCiUFqc8aQLwYZjr
NtaVsP2Fid7haCGRnjHhOOoT5OVc/lj85rlCKVuaYtFfAeraERhN1E8AUYyy+yEi
uFwQRjwuLCm9OYLSta0QqsmWYzU9TF8XOtXo7E+JdfrzBlJDZ+FEd69p8HkK70Qe
AoXkxXfocbG2u+bHiVl41Kk5F2VDpY+QHoqrkNVemFpGaDrUlzoVTTOYFrQDvnMC
3FuoDm5MrBL1KrXFImqMLstBV6I0BGLavBQX7xslasd0knG51qjCcaKwVzgu89O0
J2YMsAweLhMGeOgtAWotbldWg2ON5AO9QiUjQFCcSQy+Eajk7IUXhgiGWPsPh4Cy
pL3LMWYUJ2V3uP6oRmdcjpAt3snsJ4SHnNnqlrnTyUpGiHa69ytYO+StqhZxjXHl
qcFR4isnP63OWsZdhDmHjLSawfnhrxni2AUognpwOEuN3wG6LK0EwRSdb+fRo7Ui
ofCNgJq6cE4Taal6R7oQBOCkk+ExuoNK9wwMIsSrKYkzq9T6XT2z4ZgRBg4FE+WS
Q9NNDDVd6Joc8ARl4CyayQT+EgA1OeOv0LOvYwc/M24CV3ZDVSLwUwZOFnVHwAZj
qocHuKmnXN0uIMj27KhnmrKveXnwY5g9RLi3pSnDEIxjuiVc9ghQQjbooJw51e1I
9yraR88VpVc58tc4Lrl4qZWbhkeTd8DSVlH96PreUa3ye2nJo1KlB6ODeDStK+fP
Nl5eV/98if6Hj+I4mzkqulfS7Wwc8zAYmAbxCqfGSCQjglPiW6aG8IPqgXGAKjwy
1Zu/zi0WQC6OmdRh24hHjhB3KoA9kJ7HvkLSx7PpoSx623Es1MVmW6bAB4rPKKhq
yhgCbhVdiNKSJ3rDPUqdDNvpBMphtuNuUrDn8vJt4li+pJ7wXXA+I/GhbKV8faKp
um4e0TsMBGm8W06r2Zlk+QaxWfcIamog0yYujqwM7W68Ae04dKfwX4RaF0e3/QJb
kxPtEItlP3mq6Sbxu6uFWp2GZHqHl7ss7O2YQMePSld5PdrtEw8luoQpGkH4Ohha
0ZpvEAijDPuhqKsnpvgkJ7rNqrrXKbq8zHNVpnxjVe3Vz5RyhnwtkmSgOjGC0BBv
aAFfoeH+lrBmbz3WcKQlxgpph1GU/8vLZvJx6nnoB6uqNts6qVDB6UGQjDVMCMuq
TqshuVQYZpvruDBKyiz91lpfhqDG0XM/yin8hZQtG15F4LnOEagFP5405pACS8MK
CQriu/KmMT8F5JFB37SvxDqFDvd5QbBS/wxENpCpfAKrt/IKhMJRyIdz7mQdgaPW
RPy+castnL9A2hMOT+zXM6+WxbtmuUMIYVQ6cCLBoWt7bp5CwypvkWSUrWd/073Z
hORvZTxE+S43zWupdykN7VAoC0296xVxE+Pp/pDp9v2FZotgLpCZpCZbF1ltWjJz
xCxaWYIzCZq6qTmNsTPFOcBsu72V3S7PNhyStMgV7dy/ew942BOhPk0PGvZ7RZAK
MauwDTBV18pBxIGzI0x3j74yNy5s6ddtNzkY2G2d4zyHsGLQYgnvG3raCGjGxpSn
YUasBaPE8shS0qOH9uj/L5Fsm7A/aCnPTj6j/RrgzzJpl9HSZWP2K8aBluPzw6vS
kRwwOXKiEx0nO2HMCBjXqla7RefPRVLbprtBh5jXDW4EqMEHjMlC75teYXM4q2OT
lWn5rx/lmF4V9DRxLrrq2zPdVjkGYBCJ81K4dfxfd+vEd/lcGIc/QIaR26riBU/A
5zdkbWwNmu//JAgXq2+tAN831+64UyQgcXH2T8qN7YPEOGSRmGD72D/iGSOrvP4T
C/2OFKa/VDppySHNs7+yARnE34omKsJRTETLvxsuQnfStxMaovj+YOV4E+/bLo+r
vQOS8OuWjgSTGlyAYcr24HM24KXX66WOaeQHGyjIsd7bBMUTCTIV40A8Aq+EAcDK
KMGrWRHlllecKjgBTg+Za50rY5d7e5e71Onr87drp5fVt5FWMLWu15XT2yeNGx3f
faBDKKTRlVoFDY6quGKZy8fRTLH1n5hX66kQgKR59THJZqEnr3bylJr8C263lc6I
xn+C9QZ9ObNwNBu70jajInX0vvCNSU5+fhsmE4lwVomOhsqH7odAov4lwzeVWKfw
YgdFqzmAWHdqFBo/QNUpz/ZSHFjJC7diiC1CzEfrauC42EWv8Zvw1A2TbH6yKb3j
ApdtsfWkKsHkgRGe04bYc0P0SkWHDy3v5zw1jizUyjG/TjyLWBXzFR+JW0g0yUTl
PCkJIoe8P8Ax3BZZNh7LDlLRJpcSwhPWMUv2gZsxF0sqzzZLLSJHBj3tRbu8W3XY
aAY66QGXwmydrSwUjFnZXDM8G3OKozfWz/XeIEyF1mpET+9lccunntqamn3vQpvI
NLpon4Z1HAv0TrGuPcu+YMp0bvQYMMjPokpGDiYQKgY2XpZKaWdT0BiTM1Fg1Cel
91uhJTMXrqUnMj4NjY5+HyDdjggEpETlCHhIkBXiGvRTfqj7i0PrA3HfC/EXQdWg
y98mC+02JQpVQLWCafBlqyU0eg5TYEbF/GdEP3YM2VuxSnyaVVAqYsjOzK5ykdqx
SGHJipDsxA9Vvdhpw2/sfS/twWz2IBHKq5baWxISwwQlnvIGuH3B1vWJlxrMeuBi
m91iEVmovQewyKC9KPTvYPF/TGFkPFFayls7ExAWvdUm3it2NpphqoukmjyzUJf0
DMQekc19CoLGiuqSc4zesUxcQnJ15Jp/vN/RZh7TQ+5SD1RSM1ds7l/KfVGu4psK
ppzOFjcxvAWLT5ZwA+pzDNoSmiN29Vgy5d+bNvcq9xCDHk/9ATHoGOmvF4gxJbra
XJidP2VQnvHPXUpwILkqhfUTG0STodb0vG8sbrekOW9FJy94cLHzRMrbbt5GWxHJ
r6ewCvRKIJKnzaOQF8hDnapc89NCncjWQzOHVX3g3DL3HGduthybvYhcQwOyD1rN
ujPTZ5I/IbHDFlrOzmRCn6icxfh8e2rgl3bR5B0NWVvkMtneG+okzuw6+ChT+UrM
92OjgvxSgYPAbFGK8srO0heo5lq1LaMUB0nk6teVVS1LoCYbDrPPDR96tDfiNYpJ
+qcGELPzwsYvKHN/wsnXupRcXXcaeioa35UCRraOzXYAp9CAt+vh63Mb2J2R5JBW
9qug3ElhmzPU203BuloWQiz9Jd3WjHfNFqMjRfuzx1IRbzjK+A10AE3wBycSStiD
jTN6tkETu5geqSS/boPkNiicX2YSzt+/LIZi90hppEpfx+4sWekkRUIQRDSZrmYw
AgVyrvuIdS78F3pAweih0iYskmeGJE/V1LtP3Fo7C+1OvW6xv7E59buCAV3cFyaD
iHCTWoQpeawL49GTr4wBRbNhZ019+aIbSKHb7GSIC4HXupdcJcScb416316vF6zi
uK/L1MzJpkdBkNCZP/FVuL5eRQ7Yrc1802FS7C0SA/nhvvT0F6EQlBNkBlHVBF0U
6fZnbNEb7mAcMBou5loeMXmaAANgjkcvsXzL8hQc8etRQwWekPGNMOCteOE0xJ7L
T2QWsx2+j7MQYEGuJ0EnyvX9BAfFUaqxadm9JyFoZ22jy4IbJLE088lT97zwICe7
T2JPSJdtLzriHXpG7MJWFtjZ/ElSb9Y+FIBGhjBJWVORvUQ9yMuml1KJAKvw16rb
au7ds0wQCBk6+K94ESCG8hOHuVXwcsSYdrCMXUiQ6fheJ2qebkSvE/OPL4pOe+uj
6KFmN+bBOR8xLY3h5g6NFHH3NZJcUoTQLcFKusNL6BpAV/F6jv5PYBi76itkSNa6
RqE2vsz86WdaA3fv5k3JyONT7M2JZ116cH8Rqaw4AzTYZcpC2tjrYdLwOA3brAR6
lRCHtUho+a9W0ldQsYOwXes/MfiWJyjzSemv0ra56wa7k5HxaRaWq0sdSt7IihbS
EGudLiK1FJ2fMcUBneW6T70pukRJ1mdRmHKMesEKdJNa6l9Rxqu+/oKFO1lOtXJq
+S6+Hiz7WXJ8ZHuM12781CHYEzttWRhZ69FcrCa+mMXR5VZD5h7HKp/PkdNNPFuO
ydTGtvxWu5HfHh8GGtrrhZ4vdC/dMuNMkqHSDTt6xK4yO1KM8vZBFZvBBrDkwwCK
pWbIag978t0x6BIlAormHTMIO4rQwfvDKRbVTKOnpNPobWHWTsSyyw7XbZ6LiMkO
xc5CVSQwHyPuBuE+U1yB2K+mgRFtPMEj1Wr8RZm/emfQyQg1fEhdHWKA5RLZ4cp3
fcgoNzunm3jm1qRopEON97AuTOY58nnG1lh37O815ltee8plNDPeo4BbA6iHDxQY
`pragma protect end_protected
