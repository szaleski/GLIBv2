// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:51 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
k2+NcDyo4MdaAEgiLiSfV1uFpbhPBFlzezizO/+I3enIkgEaNnxfFA+/NOOXtH+t
WxjHYGGSSlFC6u0DRztZOFZY/nqm8T93VxNUs9pHWDMfsY7VYrcIRTWaCojyRpiU
X3Z6UQ+eDfqCR7Io0LyPw1/BkDGmIwuIVZUe2cRzNMc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7984)
nA6jIIQah+4sT04nFj8fxV8SNM1h8NR10CTInxqNOstmxWu7UJvWfbZ3G02GvFs6
jOeTyQlae2Ff7uiaTzdgwQBM608G/WTH+WQbEeb729+7zQZHNwPuER5WwxLqXliC
Mt6mkaM98fvbN2p40I5EDlz1ppOT1m5KMJ95udtL7VF/x58TRhiIfAAK9qzGxGdj
GGsrv70ifGYMb05BW/1GKEQVRd3vU2HmDfQiLJwPpYywqSq819vSeIxZmCHcG7bv
EOaG04TKCX44RsqscEyzbY/jlRkm8lti4g9HZj6PY4AN7ycgUIDC5/ywz5jr5cgp
56BGJJ8ckl5CtkPyVzrlnsVBvMbRocUGA1dU7zfroBZNSBooTsxZcH4lzlnfRyDD
4fi7IFBMt3DPlXJ/qDPRkvNpKcEARAbpmfdDsiybCahXhevcBBNcgvNouXWr2ew6
gLaLRyZKqiNnITqOGWTZf8V0gprYV3dWzKOreilYnT8UcAt+GeVlE30ar8uqapnz
acASejW68Dy39qgEH1lcLVCTJBfc4YVwIbgPLL3vHeAFEk0E9F/sOHu/Mb20W7P2
qKy+M0qAWrf7cPJI/Wc1XBPL3WUKax6feN0jY6unbyRwkJo5/kf7rg3niHEEMOid
VeHEzsgeqWj636xAs1NVu4xRvTlHUCMlNOPPw9fBvaBIlBOFi/xx3Ip01zhMUklk
YiCFCBNimbFIkL1hzi3te66GKZnEUFvV0KwfiIzcmcXgEHE2BUKefr8wyC41KCNr
LzRZ0KjhuRut7iXLnuBdpkb3OUx0y9hG1YIwSgTC4KEAknXnrg3VGmV3coqJ9F2L
Kn1fTpWCh1ZEjznMFBAHs/MRlpHF+VUBPxxCfkzJ/VC2fr4cXQPfP+6xoWUQzG3B
nsmBrhqpJOdv0ZE2PmAVgPTh1b2c/IyT+Riffkg0NcbZtMPO9cOR0uril1B5T2CE
ZURttUVEnzBPtHRHCwhjqYHJOclipy0UK6opyQ3X1vaLfIp7HFGfhXL17at/qnSr
9YZgqExQ4exa38OLUi2uNylIX4rV1uBuDSJEGUoe5F6MZaDPxVcANTzRfynnmg11
pf+w8YJXYonkXWGSm7Eks9mq7acATx1le9JqLFdnR9tvdiuygQvutKA9csNKquQM
mgS/Q60NnvtEaP91RHyDjRPInqwlp/svqOIKIfCFPJhVFq6BfFqEEmxs/lAJOL/z
bUY4DLpWsB3SyUvptR7xnLQq7hvePeHVhuJkz17VjwfpfyXdGPo9ppcJJ2nucdtK
kZujPebOgjVILN7Rftsi5LmMBBVlfd3WjtDBhOyVmNU/57YzjVmQRJdYN/q5Zcu/
4cyLLoAA+zSbf+WX0cqbzT01sa4rClX9Sl2m8HZWa/s9LNi5zJNn9ZGNk/t74eYf
AuYwI+GIY27rV77X0F28bqSBRFb6VgzBZUUjmJsgWYUZ/fWdanBnNCeirNrX+wXj
QmnTg/iiqPsoO4MWAn3jurSTgXh95MLkOYBPn2W79DdASztTU4DQe9zSKV3vBec2
MRpQdcgr/q+icxflK7K/kWDSiPeth2W+ibzrp+xqfQuitKXLfZLw6dm0lLBJv0OQ
D3HcwJAverWAEilOgrq3cp10Jk57nKxK0dxtiK3JwTXve79Q26m6zlLTqKikWjxG
dLbxPOGW7E/V5RsCCiwCl4+mfoRaQhnS6wm4cONRjOGUPQG/cnhvl5T8hwAuSjM+
5eQTxkBGagpJV+JdIGZeczf0JehEJcZZMDY+wDgjXPHMvhXBMXab+sJ07R7+I1p2
8no/a2RQ/5MVwZ7xpXtha4dLQ2z4mTYbqZLx2E7teSpSogDA959QC9M9bleO02mn
Ndk5mKe9EQajCJZe1J9U2CcMk4S0W2fmQJBBWhXdNgghz8MTkI/X44ySbkYKJiRe
TF7cvxL2Y3RmBHLsIri8rW96d21GVX18GXMGD1CtEw+mFg80TB648u4coodbkawr
x9maBlu8ErPv3duzNLWNO54xCMQ8DoUBHaicSsK+nJpfrPv5y+vnfsyT9sMr86ag
A+noXyXI/5hv7i8j1TdeSaNEsXnIYpNnR9jtg5U9AQpjzLiSB9bshU0d/EVf2vbP
EFTU3CcAW9PvEgotjCR1767p9YcMqIhRV+lcEkGI6yCnKfCcbAEku3gTF2WcE7xw
qw+C0q7lGaDIhZmuh8Lhi0V9C+LxLH188RW530dMFAT8u1/rkO3QYRkzwsLtQ6vS
pPiFNj5fqgt6bxrUO2VZr36g6afzSrsrFEra5Sb8TuDTYEk3zmjoWg8N/Ok+CMYU
joTFQKySLkSCXvCZ0pYvnmCEMLbqpAifQwveGBJkl6ANYVQA6cJnboEl4ZbZL+0d
eZyqf1JnvXW/Rrm+rIAn/xVIXbiQk4cGnCuNcltZgzQGYR5u1EUEb/40x0tbLCcZ
p+EQhcSRnQt3k2VJDdtXB8WMrIthAM3MMTSRFidBwqkeFQ+TeDQewsvJ6VFUbBoR
pG7NKWL/H2tRfth6PkAiHKNiJyBcFnFKSycesbpqP0WmzWTmmocVZDJy6YHoE9UL
iFP9KLbo+dOMbtbVeKq4u4mn6IQy5dT21Q2JinZzmDQDvk6vlwudiTzHpJDvVKAG
UwixNRIO54fWpm+mY7gsUJ20VAJuiYVEwBZJHy9Ocf3dkkRNDXbeypTI7BlB30FZ
D9yeZH2HSHOuOw8vY4cheo9hL4/cHrP6X+YyHhU1nocIZENJG4y1rsdkp+gmdlg7
b641dAOxRTiKm6Bpb/0LamExJvD/xkLw9bG35SPIfhyQwzKIimiuJLzH8ls7YTkn
IHfj50TYxshTZ5XsJGNyG/vWNZAtrHLvd4jdqrjaKiHRGn/J2EbzODlA+pydw7l6
vn0P6oNWtlm1JrhSzo+T//C+6mLhzUMSx0Yhwh6GXRMYgVqR2y8bVE/GT9TxSoxH
eJYvLT2CamHRzjtFZDMc87UJ7+fe0XZvgFsLrb5WtccWDhEvdqx9XQrdEKyJDCD6
bNIUwQd3/h2rMhoExkHr1x69s9pvVZ2m3QAD6sHXTlAQNbZpLrQ3v5oFenKr2yDx
g5r4pw5nwYoPgct0R8Y7pUF4ERJ+cDw+J0Aru5LLMyPdyDIE96Aa9kiCqE8r+2Zs
fXnoGnoovQx7fJB4HHL43i7bNmlZAwMfTN/bnneeI2qKK0RCk/pmhMW6KvcQwPDm
yKaD/PsTImo6XWhbtpeU/HMuWMcBJX6rPuBHuktkkVUbdTiij5aDK5xWIDphOSAy
cyR9LLqciNqFmwiOCLpRz7TAY9m4T0ZMQdicmxpa0wQBHZGN+2ebWAixD4ynETCy
R/5R8EEu1Oj4yctVDOnQMbOSjeX0WO9658Emld2ntCVE470Qis3Y3PfWvORWG2/k
/plYb6ia1CBOXW/3EId2IJjE2auCnWLsShKiT9QbqgQdGm8umzkspPpjtCUXWQ7Y
RXEhks3wRNK1FC5NxYNs3DvARpvhMS6Kv4lt31SsrWuirKBUvJ4X5jjxTLqnlkBT
CTIuQIBryAI3mE+dYswcf6WLe4UTY9tunFtdZDSBmfVTmGVoFqZROb1rUqmbpBzW
JSps41XFFmLADu1oIl5AOpu++2itRRGg33CGaZTbhn/Y/ytEKQ5UNU8TTWhHzyMt
QJI6Xkyj9bJKIw3XyuclPqfFVD/Q1WoA0I31f9YvEIINLEPO7w5UgGtnmoAsGn9s
9T20jJ3lOBUOqJfJ0DysqcblIl7y2ZkdkMwSNCzGt7tLi1G9UThJpLOf16OT99rH
2rceAtG22bqkyz9EhZiIFwiU0ixTE6G/AipqRleKy2/y89kHEX03nO+3/+kc6ty8
Omys6nWZzpWPe7dGTy2/F8FH+lz9zF03JUEzeJsues12Kz0tsBEyk4FLojZLoQ+Q
ioOLCfLrgVhTlI+1OTJ4KcLUTlJNOf8VFD7Pvo5q05tbiiQoIL/QOvZWd+yE9z3W
n87MZHEB14RFIvJ8bXqDXQvzOdgAtpYZOr++4VYzGfFmZnpjHP7Nmvdmn4ORgX3W
CDWO65UTuOBImfYtJwZfNv5IwObT6N4CeMr9sl8HQuzNaTrow4Rwh8w65BtpLJds
jp6L8mUDc0iuThB3mCBLR4F2IiD7kUF3A1dHHepXF1RbBNld2kQue5IH64jYKicY
cXtB4i6JsYv7u4M35afijpptxZxU59t+RdkRFZGPeEXMN3dOE2vKBh77yomkOg17
0rdQuhYDJJOj981Z+EiIx3ddBTfKa+VYcOVuc/xGKOI8DZ9J1RWDInIfXV8Y2lhD
ov1mSbZhm8LmTHg+3gVSByOgt4+m2Bb46jsjCkYI5JLSy5DgHze8EjRbUh6Q7sTB
VIGOSqklopCuGXBsBF9AnFLCA9kmWrlG77H6HsKQugHVDTcu+WwU+vpptdsiD+Ku
XdtGPzqn6UZLyrbPlwwIskVJhKwOBjfKbmMItMJFXnrpJKkmbwliby3952Qzx0kC
iFAVQ1qByrv/X58WvSQWckJ13eHYlGvz1TYHDMcghZpU038/kjMbZWKxX//4BKQj
gOmdv5VKvvRL/SvFX9QKuoi9MmG33yaC2FtvQ8ggKgpqLa8A2GdwU5bciDXIQPsu
himygngyV5UjqTai/OWkCoaBAXsJygjBCwii89rimcHLkOTFunr1DsIAvzn8Gc7S
D1Y9JGzoikKc5fQr/61bjuct3edrc6ixkKJeiJnX2CWqT4U78JIsyo1l26XXA3K/
Rd0QBkYyJQLYHB8T7JeKBGkQQvSjwc45MgJbZyxnR1OPvLrKvA1O+aHPDt8sHgXZ
7C251U4UeEKP4lFe1ghJt22Lx2a9ITpKues88WOKEGhULla/UfR+rSbMPr6NTS/9
D6kA9XxTWAr3kxU6R7zIQHEJ6pKnkNpby618KDIpstZcnOgWmTskV3q0JVWm7Vcc
B7uRMeHQvfyw6yNp/ov+FozVraffkpLYSgf8WdrsmxtBKrRoBGOqFIE3ZSNqO0ld
FZsM1UVCpHbBYIZWoAlAMB/fHtLG8oq+19RLG9rena0vD1a1UIihlrokGazUH3T9
v9H4zog/nONADpWF8neFO9Lu5ACRvlSGUkuEXz6cu6BD6Eo/uI2wEuJnDi9kb/sx
7ccRypWo24ijV26MkFCoabFtQyr4+kRFZJe/qjKf7LwqCrnv8+IQt948rX3tTM1W
G3bUfgek2RGjTy3c2dfCMNdFLUbQiCSlHAiIpZLFDl/Upl1oOd0H68bczv/yrWKY
7s3CXbqJogDtGwVY7PZiUJABUlGS9MlgsWSAwVG+M+bZBKerMb6eUqQCa5l1CuSa
DQbu4k/iop+nMuhLK085yCtw04omJeLQGtuYFAnJCMKMs3dkhR9bSht21+oFI2PJ
9vPwADqtywNRF4Yjcb3AEsFFXc2UrQlXIvxNLL8Q1GS1A/lJNP+d+yeWnQGqHGmZ
SS+hW4WrPyAuFWfFUXRpe1xJ4c+xBbCbh1Fq1pqirE62EjHtdTNB0Q7R1CJ4XBur
3vfgLeJvdgANANY6OQ9MMrI1+fbQ7LIOm74TJtOky76s92kRiQ0Hdc5+qe1ixiJ4
YX7wdAH7MtxFwbw4Htuu2YT7zbFL0QkI66aRuCPZutHsfp6wobNvxRTDYXXHxBj2
0lLGqESG0yhidHS3SM0z0OXn3FWmW2o/LOhF1UlElyffpmx/1AlgSFuBNcKp6L4h
la3WUsHq3gYGhJtgq2hviMKOfnPw4QCD0Qrmj3v2jTGXgQxo5jN1IlUE1AuQ5JrB
MwzNVyylei1pjqaWDkVfHqz+9L3vhtFrPQCgYB5T9x560N037ecvHTP93KPRrDEe
cqYjJqeAlH0oy9HtmPyUhoukmV/zeKTVhxfpFMYEJfQTS5pawy629VkRsP21YlS5
LtnFEHbRKRjocfZKEiUbY1wNt8xwi3A8yx8LnowA3ttUnkDQ2GRavoISyN4CZFGG
2jF7+eU5L/iigQxx47cufjJuz0ftERcbLKSZabGiKBGUGXGqHt7BcbrMMwVQX3oE
nKJhH/ZhIOahuN291kjWSQAAcEloLXdU4ub2g/q4mblp7bgAz1gERT8PGM/wr4sT
LM2TaL0gXB4n1dmNEYyygfJfc3xFZCaXy6oNbhvTZvGTd6MuwlPF0jXltgnXcQEN
ymWFU2pTr3GTYxeiSCrvVjcFflQozdzrt+LtldaVUaa8E7Y2cj2mT8Z8rgX1PJ2X
nQAY8anjr1DZRRdSQfTvpK4IIeLhRTlP4Fa9JwkGZxJ0RqwMEQhDJcjKEM3OTrj8
7iniGNzuPJheFui2PxchMhQsVlNE/homeAiumRxukMKigJsF4XOBYnZiuVZgEukN
tunPGoKJ2x2P/fjwsYIKQYNBNzuFRvajKXxUJvkBipjoNCbbw/p7PcLPLjtKyPHE
REEQtrclLT8yJRpljykyYVf+VSMhfPEYa1ibMCCdtgiTPDD3Or9zthgEtOHh4PLa
hnAVIgE3Ax4oxcYrVAYuHcWnct9a+qyB8hl2rBMUcVeItoihRLTKN0ItRBrQPCf3
Qxn0+WMn/RQjEo9aXtYO5SuhzoB416/DIxa/15cmA/4okjNEEE4QLShgbd3cd5kP
+gjlnfIqXjdzjcOBubuMqoYbfvDev0b38u6AxBTZ8cMhm3D4alzGfYrkcq5TXnQ1
yb7JJeMROX+m8i9G6t8lvY8bX/140AIr8mbbaYoiOmY3/7gOHfQUNj0HENhH+xoE
ku0vVLfU9ByODIjrA32JQ66uUYBVNuOgQRumZynZ+BIVR9oC34oObcidjDkrdd5f
RJVaEZz5cIPu7RZWCEPj6WxcJf56fMJqPfyBJSIp0eTgttFGqvMZI4NfQ4AZQps6
iix7BXLhya6bmUZvZvSDU1WsfXN+6ysU0axU7x6iRMbYWliMHpAQ8goncZmoSFcd
SHXy7UNusz12UhvIEIJw6DwbJrIB0g+L4OzhslcV2Y3mpDrpOZH429o6B9st0/Ip
oNIPNwLh9XfPXDq4Dl5BL6gz8DOpopNTloaWfjEAutWeZhYQTLL7hmxQ7Y4BUzh+
hbAIMHW8RQf50EG8+K6B9jvG4ubNkCm35C9s8PbUEPnhg85Asum31mu/II3Jgqur
I6m2sSBRW2g9dLKt70+RR6lWQ3McElyAnBptFWinrszwRub9052wxk1a6xcZbnyf
oWcLsLD7f+h8lIZp0Y1ZxNZsxPVpjCFIbPGcfFptK+4JQrCnaGmBmnMasrWlAYyx
zSZdEtplOL9xJxGz5Ky6Zn1gxGECO2eu3XthHe8xq0vAHdfwRK2KH/3bumK9iKbE
cK7v5CXWK0KgrqNaeMksuY+V/xzHUDVRAcls6IX5WZwiMFJPNqedsMdBmHjuPpsX
l+WUPf+Boy9mPn6JyBcTJfj2t2dl2JkzEeI6c02ALLODivnH3MDwhrRyVNEl5IET
JnABxhYyVhaqB0jP2NGKwOriwfH2FEj8DIhQalNZ6qIJ5Ty7VCRsdZo05DzSjUPa
IYxMK3BNgS7HG1zm+5wVA17ATmwiiw3mgwd9CbckiWnfHXpUysGfLr/y9oKhjpMM
DWuLpRGNHKrEbO4vPWtCnSDTESXo4Uh0KhrRqUeJZsPei2Gnq68cCDhlMhRmigg7
RbfL35a+BG9hmqBKdb4jzPGYKLILV5wHpmXHcGK5WYeWiVOwSFNBLLmUP52RpZiY
sm5O9g2Vbn1XR42HjZr1v74WisbWilx5hK0XTV8iFcVW81y8T/Mb0P7yU6bjRXCj
J3jZEf5FZvuWkCEF9qcB42H0MA4Q9NRhp9WloPBMqMWUdqstnwuvaTsW5ndHtpMc
D/R/FzYcIs0A7E42E6YLVIp3/vn5v0VjQrljEqvNuSvuFHQNP+fv3zHP6po8OGH0
mQhR3+4Y/YC3Sk+vL/UiWT0X/KbwGRsS0RcRfhmzLQcrnnyyCl1IfAWdZ+ckye6q
BvzOXX51xMihj7azJO6Ahzmu21t9g9fzvTb5I9bX1N2Zu8IdLj1RorELllSwSCnK
KRiER5BDijw90H36XXuKpvUiV2Xv1u3z+PCm99WSf+Na+itI0dBPPf1cDRNuUwv7
su7f1uPq945FkelibGPuWLng2eDjaxHfGPLcz0Vr9JvMbVHTb/fiOnbj+Ituj/sM
8pUNa+K+6zckmZZDzEDDxTLyPNFVQpB8A+OzxFXn/DCOvWNbB8dGaZSgibDOoRNV
GcLBbUmBm2LCIWyAQFmfOV9M4nzweI0qdNxVtROFLvePIYdjPJAiAZrRHlaWiu9f
9TXrscOK6QHU3rJzVCd82D2RnekVst36fAi/8YXYDmdzJffwkvFLyYagy981ceI3
REucYlHQ/DoIvUKipxRNn117JSRXUmtYNMZZibk7xXoLb65hKgm2W/lxMMtwqznP
hIgnwbjUAIjamHVKoDqRZzJDXUn22IRIbZwiP1qQcl6Z/pUtmT62OWvYI9KUpKAU
1AvJbN/GUqbNh6v7gAMvJ3wZf5JWBtGN2ONsRkbSP/UFxlxEhHRdFTcYTW2GITNd
PTgXr5Io+vFKjM6TPkNC9p06xr3VaQktd0MV0uVsytw2quhBigQ17g9vqjxYSizq
RT85kbqOEEz9Odhi3QZ66DBSEjRHMMupkOWjdCQKyDk4ZBCo2PFKgqsc/UsmACvl
tQrbSsl4xgoxGR/FA9I6ndlMU/xYfCoV7lzYQHRwa/LqHPq2HD6dJEEPlKGzlb01
4z64JTYl9cmnNb8kztB76IBEvBKbzPRTiEYuIWbT9MfZNQIMEwGG0g4JL2gOh72+
17xO6tK+CtsHXPEe5gNeYz5ZZX9Um62HV2NXJ8V6sM87kEWlxp0i+7DHyUZLpstE
wt8TiRDCyDsaNMRaZQmv8qPcc5gyVbTDzsu2u8l+SFQ59Qdr0MPQDjxHHbIck4XY
jKtUlLfQNKp2tyxhFvHkbL0uBzaVb6DdQti5foWXWEnz+5uQXe10GB9nauDmSXIA
xfCyxy0xoTH0fWwtHUdHf9L52of+0O78SGJHgKNZVyfVbbw1ZS3DloZkyKzWSBhq
8m8TfP7c8ZbGRCewmdrwsTHnjpba7MOKA3t2GOkaq2MFmpWuUydpTbMF3ITX234G
hrmXwDAzXIYhWk8oJeOz3rzEQwMZ4TiptSV0nV5jXDYBcqkqm+yx1qHxzRaCu+HH
jnQpSvN7NgY7KY4vVJD4ycAknxgxUBiCmZaEAiVHAsoHW+gM665LZ2lVQqjYkhFF
3Kl8jllyZrDTCChx0YNvXMI9440c58n59ux4KnWTNTZlcarUw0LG89mQFaSdOKG6
qmR61NDXz/KDAh0tC123MziT96D3WNOEPEodWDQLuuSKmVz+zwxs1Ex3cpUFGWI5
mfJNbrPPjPhV1QbvEvo5nZcwbBixDLTJ5cHxCcw7xcC5xZa7yKwIX6vf+XFm5c8e
AGpVJWVzFFFjgd5cJbWDdPCHAk+Cm5oJMs8sDeb8Iki61QMeilB+cSibWAnm4sVG
8e+1yE1WyqUaFXt45z0BT0v2/FQuyECGKcgazQNTR01XHw6ZoVGsv+oeglDrPAJA
A2CwaSRXBpV20v3bAJ/hrcTNLKe1U19LK9/uEaIwxmxDzR+Ioe1iKfqPcO4yKDTr
nnMy4uR9MvY3XWhF/SzUpuUjm6SGiWpsJJcIXquB7z+qUPBIPdtU9GQIH0OH9ZZD
G9zQL6mw1I0nABIEw4acaAh3wD1fJ6Sdi5+v88RiMyQLk8aUKFJV0Z7h3ExflKT4
LGKiRb1RrsRJFdWbuj+YQK+s4MkodquPKOWdgzUlllkTXXfwJZ9yMwvwckP5YzIQ
K39/5C2N7fNWYm/aa9PIP0lXWtTfuTbgT4Z4Juvz0oGndlen9xQS001aG4VrNPOg
WDWApAg1O3WXP5d1ToH5Rp1ZN/qlikA8KNfD0IRf5HwtNDoPp3tlyq+smVzdN9Gg
u9BEQCne11RzmztvlCB1PzW91H4UGQgxv0SbA2ksRET4omUntIx19g3GmaQ65cfn
jvmYNgbquy5dDU4tdcNx0Rzzf66xnpCJWIC+cy3Mt+JhBQehSl8S595ln+5axTlI
30YtaqKh64Jq9ZbLA6cNB4YfFAd4oSGA96B2lx84rSlDZYhf0fQDfeY2NCy+0ksO
yo3NGDekFql1HmYWr1KhM8SIc4AVlNupJb/J1EBehMODi0d/2TJVCIwhxaUaoXnG
eH99rQCQK/LaFGa2e2KClWiUWP/n8TWLtA+dZmZPHLlPjIDqIXWICPCF4QLkg41Q
3C1FJAt17kzPY2hmLiBIO2qsmkmPCntfiGDB9TNKR967qa0iAY6nfBuFIPMScqVp
RqSlSjhwIyUb9+VstxcPuNXU61kMfVCkPOpTQ9a2B7932DBiPK6tdUg3sNnfbzGx
V+Goej/z0D6r7ElqjSnhxD5o69vUoUGglqq62srmF5J6IIMhhnbe3gXYvf0dUZN1
mrPogZkVeGXICtMjL0UsjZI+mSL3Vh7ZvZzHDbKFZLaB/Olgixou4f79OxT5tWPE
2+dAPisV/zzNwEf26XsMK+Eusv617poarw5v5QBKDn/qwXJt87l+h/V6hC9biZ6h
mZ9UdsYw6iEH4yzGg5v4OXs4fu4MkB42yMYmAtIJ7bsQL+OPJjjAHk4AFojA5gwr
xM4TCCOujeDrH5AkxPZVVg==
`pragma protect end_protected
