// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:48 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
NwkDTzUqUuctUnZfAQ3E0sdNSbPuyNU7wNkQKvuGZhqis6sYP1mRlyVtMsaziQoO
XO1TN2FfR/+XUrHzhYUNJHyvGpTMVfGQJiTdDFJHQGtCLmN8AZaa+W17JkYu6RdG
0IVsEuEb2v3tFgu8FEP/FTjbs7urGgkymUspRvPjSAA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 14016)
1TW4K+UBpq8SpmDuopMl2sngz/h1fACHNInKyHlG9BZWjVhqhcsYbek55s+BOgEx
fMPMhn7g/S+iAaOuq7tn0wO9mRHuH3+Is38+JPxx+PRiprez4xoQM/aJBS0P4spv
eamQL8AYQRbRA7AVGBc1xfFjbyq1KAOGiI9qQbdSQP9IdTrfgmV6+zkZJU7jOMLp
hTV/hOfxaHQvKN2j6vMpTL/5bAkCFcYxDzmn3t1L5l6UnJuLweMVgNrLP57o1Zgz
4m4aI+OJxVlKzRveXySg5Evy9dEwaj+tKW7v+dcNsMb0RZbgH4WLLoKxmS/WgknD
7xgcexdw0YJftUNjo49uPHRL3cxNdGrsXqGrY1wnM1m1B4P6b20k7RSmU/PNfTOk
FpRQ3VcpAbwKX0FH8ShNluHIYBFHXUFykttbj2hHSic4QaP77kPnnm/VVJPnuOwC
a+WmBO3TPPbVR+VrgbXdnieJtu9ZTkAuHgaLQFD5H3zqOaj2zfF0AttGvR0CFvHd
2KWLfc+glv1/hYIAgczQ10eQrVM3IP7SeHXJM7mLrxndLjfXxwC+ue0c5hmX2Z0b
1ZMg5gmb/SUi9IVy65iLvSJXIxHgWmvF9E4IRg20ll52pKn+fLxS1fNxX1bld4EY
zOKC/jS2ugXbutZyDn68W3ztInPgLl3fbupiNAJA6cq5KngUpYPyd05wT7ARqZEF
hr2vpo1+TsfDOxE/sS2bryAbyHLbbuATm8rF5az8PHekBR6bqNv8XCT3JnRBfmDY
sjv4e9bEGl6QTVvfVGBfaVO7xWYKKNuBAlW/LfG841AZ2z6S6qOG7U3qmM5L2Qlc
hBdHx4t7CvYdOnP7obV4mQB18/FsvkG0X8oyyDWoOgDGyta1Llts2asIVa0HucJh
nhNwtxaJE5PkwGejhtyTvr+FbGPo93qVjaPZtMgaS6YnMzKJF8qS4FG8sXR3XV06
wUmssNzG45+L5U1GYKU/aNqZdCV1TAgpMkjPH2DbmZXtBC1cCWkPRfVPoTskqion
vT86KfdqkprQib+1bbL3FpGy/zCWkXgwvwU7S7a06fEzHgj/cnCeY6K6JMrcgShL
h6yb2WP71G01moOrf3Kceh+3PR9xCfsPAP82+xGJHM1une1g/8bAj8pF8L0RIPSH
RXItLc1N9CzinOKgLejRewAkyXuheEl52dmJDobHqV5gPi4hE634HmKRbMEWWhkg
5I7tH7jUr8i4xIOny149kaurXWd7K+HPi0ttHRA666vYP4B/SURaf7HlZDSLe3Vv
KC8aYcoXX2LjmNCy3PiD9M7mIfVsoaiinl1QzwuzbPCXpn8DHjdxQJyX6LeFkhOl
UwtkzpTNd99JiA1MJsoEyLDr8h9nPPXtgvLWBwAI5m6jqqbLWHRA6Ob7NC5NaxI2
E0SFfi7YxF8FXWbm0s1qH30/WA0jjM27b9J2pP9ouQBP35i6wqMLO9o+zCvf7PI2
3gzeWTYaPKM9tXjNEj3BVAPgeI4y8FCB2dFBPHVoBHnuvarOzP997cFeB/r5iB17
iKHSkKe0y4oL23Xc/igDjYjzImLp6eW+Tjc90aSANAoOxwgR6P5Of9SKC9pdBVUY
CMLTIaNvnJkJgxj4dSNuV/VqeOoZHcqp4+Ymqgrkbrv/zxrKFOq4gq5xerjJck/e
7mCEYU+FGI7IiwxW2kzPjibIY3EKQ8DYaQcfHOJfhDSjEJWNzFl+DHDUJx8a+giN
43Deip9CCIHzbwitLwDljP6o5P2yl+eh3+hY7s80xrVof3TPtVtJIZDcLSycPzfz
n8veo4t/JzhJpuQ6UcQeT0B9DLXDZSavgaGHG4yZHOb02fVd9h3JP8Xu2DH1xJmi
xCIDCI/oDFhNCGiDQRfAIqczgx0ROlQhszjXcDv7PVYkPPTEJAGcviyuKEnralhC
HprUw5ehkPqQa/8CmJ8b4aPeaz0d6H59/FLQja32hSoCfbXD9JPI3KpOb9C9relJ
OAMEDBobjMGQxPtb54axe5yNwvZvlvNkj6/Nnb8s/36R7SeCzJbq6dDawp25xMRR
4qDYcPZipy4af5NJC+l0i7jmJwT8p04JVk6BOgAJnxO3ut0Yst9D0CPNdwoxxY8Z
+JF3U6SPFF4S17xDwBqqzKqn75hzwjDuxB7VPKqGwhr5RY6KkD5cMofe47hemBRx
NEFnduJnL9NhyIIaHGk7lt30j9S1D7VpHZgVn/N3M0lNCQkGWr8f3dt/v88utY56
RJKNU/vc9nE/S77zjAjlUIlxgdPhbNnvkq53NLtfrol9JwdVQfQha3lri8Cl61N6
SWohKI/QpBIkHQWX8fgi5UbeCbx4NK8uEzPiShwKfDeXBPcBhGvGJgQfGDZ1QyCz
ma/ez+Xe1XSA8bqzIGIi6R8VFxKXMPzbZA6pulpsUhCR6Ekf9FQXS3UprNHFFN4H
Qiruan3t6PJfJLQjd6gTq4+VnpUJNcCEyRHJ4rfbaWCyb6Cb+PEmfmDvdH3JnFwY
XDCa6kh+m5exoId7KZD47SpvuqwEwcAIpaE+VBcPPCOu5ls/7AOCV+Pp4RV4hoBP
K4O/byAem44L3/A9ZjRVSzG3mJvkFiDwua8nPASd36p+Asz0F8zeHJYRgKvaYiA9
2VoqNBQVcIeA2iyJByIO5ZAuRCy6gOPtRr80W+XKFHaEs2jPrDLisSqsyRhZmLuD
dxxQwepyMCTv/cgFAWxlxCw68aH+gKGdDhN4tdBnSJanbREjWgYa1g56k4abKsPp
dco4iqKTrMkHt5II+w8dlShn4P3j9SaKiKxtiJCcfTS0hECqf4M3wjjbazfGKXge
TYxfINPHFLSWSW3ErY4pBxxmOGlS0gDH77xeZKJfoiSlCbjXPRBOD3hg91caZsfp
jnpcQEktVHkXJIg2W6Sg8w+C4VuWAKrgPG4PMLtuYx+Yma4yLKE6PN9egJrqJJY7
V3F850FwsJ1Q7EWlO7s17aEg3t7AQdMa2hTlsLWbLrtS/7PyW2mVtJUaCsudrXKP
821bd6e+N9xwW8Ncy7ugBWO9eVxL2bZWwuOkwwZZnRltPZcXWEcafBBULvLobG4F
sa76kSYT093weF3kmx4G7erof08+RvgCBpQaC5zrGOmvGBpIU556qs0cZ8sJLGZg
ShhIObTjuvbXy4VHFJ9vNIOxJxH1ygefK0T9+N+ZILwnxfx27Teu/nJX70UQnEGd
T0oBDodh8ASNGD/2cnPhsGbZicl8f0uJzpABMeFsiir8aZqZ3qCsLLTFzKItAbDp
QU12FNreDSmxx+OOv0HgNxxyoT/5K+XRlPO0jMq/a1LV0196iqWaR0zjtCeHX9KO
L84Hnmtm0wiYV8/bTkVPnVRECHw6CWAEe4znF3TJ6aGM4EGoMOvgl/X/Wh0/bzM6
wZRQeH/zNWAoeCIG3/V630hnnyzzOViilRdFR0ZZzRjXbijijlB70AEF7scvaHrO
6mRCDkeefWHG7LXbRp1Xn4bnW6cdFlRLFUbTsl4H1FVRtnr3nareDfxWiKzH1SL5
HEnrlL1KbUuxHEfN35lTZhV/twOACMiev/Z2ibjCQCS6n+Xr+inbWvOjgkxsweCy
AfOKVLy3LnhxWyiyC7sTQ1uD41oXXLZZw+C4AN6BSi50tCBNTGWO6lGGrlF2DDYY
Thl43qKXaC1hE4qzDy4/9SLKWdce4717mFyeH+bWg8RC+vooQRDEL0MoZcm/xufU
dDBrm2s1QS2VI7gtvAiVBR450Yb92f/48UugsjeOHHntktsg1FoawMt4khVW9xC2
oV2u70f5IIR6mdXtxxQpsBirvMQH/dLSxCcHC8Iu3vVIY4cBH9apAQkjKhTAE7GO
B9c+qD3afRr0aywXTl92+XCKk19VPSKZAKU5mY7LeKMYEjZgWKrdEg+3AwY/JUFZ
4Km66+sylzmI7bHHGRicnVbXEaDhpmcJYfcTD1stvVJSKM35wNcomdmlxfYsaHY9
GeMcRjAaM3QGS5Os2oB/W42XBvpk2ikIA6WJ/yIe0akyUzzhi9iwTase45jkhRGt
vzdUeI5GCy/S8sIhrkD0DJwh77BsEm2SacO/W8L6hph0IVuZMsLaHutEejmAY6C8
q52JyXT6VkLX0uXUhsX/p1xARQMb2g917j5vPvsElGxQpgs0IddpxYx4HpXyvjkX
pn2RUNel/iitk/4s7dEJBzEp14UUB8ExZmGNWzELpKTwWA1uyxal9beFYxB7Grmn
7S0GXDBMzAfK9cPU6d6SAShvY/naqJz5DFvCFtntDEsrxSFZJKjCCHXQNi0q2gS0
dcL0ZKHXLP0I0a4SY43MJeh/+CXtnHESdGjzpV7rcsIZQykqhli7WZR+LqcetXcg
SruEm5d4HX6kZqNPmC0hIAeHFYMO2ZVQdxKQwC1atAmiSKzs0WUczEDDtw96DWg8
MJBQLTHYwRMNpDFVitR8GwusOsN0leER9AOlhB8a0YMAHcYtQc+Pz8VGzztRiuVa
OtZaJHyjZr9dPFvXbw4H4xfpq5FX4C/w4LwIyX2dlDwkECLB3glyXu8wB+qpw2/V
byc8wAmP7FELOIQBEYorsTOydqN/HVeUKB0pcexAy4N8+Dxmi3obukjlrJv+N4Ke
7tFheAem0Vmwtho0xSxJfl1V3qiAZ/mYs1CVvvNUbLkK+Wqc6xStL7xyjHWvns2R
Df4xU5phndTD4SyX/GkK/n95Rwm9KA5989HJSW8cRjKhlyojD81FIq6igJh0TQMp
iAZU5UQEDG99SgqkUTL/6upb+RfvgywB32llNhs5oTT0s5LjM7vFrn9jZOk8j1vh
s/Zfr5jWFNtBwdL2Z7DAtgjJINxnIWrtt2fuVa6waIBXudMnMwtgVPxxlB0Rd6s5
Vccg9aJRzfYJdXww2nEaIh5G54j+HkjlNWs8bF4Y5cChaRQ7nUZr4MHPE2IjDZ1P
9cSwcpHZrLjkkl63DylGzLrp/UL4vg4vPmYUF7RhEnGfM3EpXcDNde1M2FoG2Cp3
bpUSH/KDhF0MNZ7HedBz0hCrv47OKacjrKEd0+3GhMPr8Rn/oF9KPFz0J/5Xn0x9
lS+N3k0NqL+7nInbOJ/UgjHVl6Xlc8Q3zeGYgjXH6QxfTa1hOvxyj1t+dvuGOzYf
4QaOx9jb7hnr9q3FPh3jKWhe3MGOthXrgiA5gGELVR7X0H5rtQOny4GkwyFG9o7b
YDqrbKcTPm9s1D7muaDrSzaW5Bk1YStB+BcShH9oogtDVX4VkbnZhzJR758CJvCc
3nUs+yjSu4rvxU2WLohdVyTI5Q8J5tFPzhniQ7/qortFHfnKCe58OIGrrIBCrSde
qzJ6nzSsZG/TWgg8BUQ6wNAOA5Hn4NCzIDXQVD86OjEv6fHjmlSHPwa0DyQVUSD5
1cNhgc2PaYdoWMpn/a0dndH8iRQTpITW3qq5qkLOC+XUGzHlMCedLXKU7+lQfAFE
eMNWZmfL6gAGDiBxTccEo3VMHLEl35UT0pBw1DgCsgdI4WDDXWyRIXAhPPOW6k1B
O1zZ5/kDjoDwj235oD1kfm0MeWjz2xMJ9VI9ArL2hxeX/MfVU5yKtYNrlyx+MrPP
rhVclYsMbtPid+Z2lkDir4Gqcf491Ony9cLF8IqNcIvdODS9Jf52SnGjBim38UgX
5VMeeLLGJRpZz/zDiePZMH5hIQjXYOdnvMCWx4Xemcfz5FJmGPs1vM4gbpHU1yOK
Xl10N+AT0wjlWm6YddqeZuNWYa5MnXvEdPKgps19IcTPODZ84eYq8PbHN2EtImB3
fu6vbOOwa1uM7SCxfFtq7SHXcgmaoYlqSsvDLBofEatoedgGnnSrETZyBJoYx2dr
k2PXp+1V5QcU9pRP9H8cEMppcCHhw0LDgJ7aitkZJA29ycpEj/syStbfqZc8dGAu
EeUAt6SuQvOhQ4JfG4jSiiwWIKu76GAIBWdKQ4+niMwXyRGrCCMKQCZfuL0YgGTG
QLkOih5NFIr0DUcz8UEUCvo23zGPlZPqHCtprROaVsaMXGNToCdeR9oIeI4iph7B
wGADYYtiOEzTE6IB9GrqJUs83RDFRXpWWdcJC7wmf4ury2J7oRUodA+YtWEJ6FJC
pxBw/kxIH765yb0KZy+vHRszRGEjxpalj3RABCxt8vNIa9J4fhz8rWjN9u9dskim
EfhXl/iFz2cYy5vq+sOFccrBO/6sHeW1oruen+VoPVzGKhwZ0PzkWYcvVak/PIEM
pDgV4KJ8kfBj558EhI7d+953bkoi8tSCyTxaJtaEfRsfS5XXfsH/2llmnNlRVAMx
98cSkNOD2c8qlz89kOXv/m3xijXkBSgiX2NileRddnum8rNKdmKeOv3J0ZyTcNzv
QQ7WahM2gKwwWMj1bPUfJb9ITIOW5yuZZ3PFKL8bhkFEsB+ABHiVUCiRjvfYoy1z
BJ5K3ixB3it2Kwyj1hapNgeLK+Ww0JTOl4HW7QIsYBBdrHrETqH5fp2gnsMUkES3
WmxjxdgWsnvDvWTnh16hwpTLd2XL8A8Sy1TJ8jw9cgs/l7faUGFwdelVu1sR1vLt
TXur++/EHIk/XTXFbIOq7e+bQLq/ODyScIyjpGbvcl6hQZtEs5GtI+U8y9B5sGEG
fCmyA2spaVUenRvzyVqR3BJkYsgYHl10kjknhtMIeaVcdVUdnxpQx8wMG2zlSQzL
FdaQsWCCMN98/tuUdrZrBHpjjh+a3TuC6w1bp0wfw0GelnS6gHfGxfCnLBC3o8KE
9Zq8lO6MWJmFeTdchduz7M2lrsPELlk0C96VKlLqrRW4nBbIvpkjMDXMCbnO75Vc
3HrN04S8N/etcnKygs0xXGx5T0hW5a3y2XsUiP2UtfpZaxeFGIGp4IGYrp7/T50b
Nibi9w+uE3Fj6ovSKN7ItljxnCZdEtQb8+kS1OOqUdtRd50kUhSnytfjkChs8h+v
jOvH+NEhYKg9QZ2zjvNgt0irI+ljujg6xQM/HOWkOFRahY7KPnK+lPjcjVQNwirb
RYn4a17WA+VwGa05cOuh6+I/qJCJ0U1k2rOiiriGuj2kHYN6rPf71MxcAvZBdUrc
2FeWHAaSMxGUz20+L9sTvg8BTle2ZH5s1H1GRQTCTXdx9WEM24CSTSZV1YdyPeHG
aD7KjKDQZj7LS6owjgNkBPsCuLLSivinGN8Ym3QNPn80hyUQZn+o6729EJDzIGRP
LnkoUcdRCmQhKDd4agMIhF7vr7fjvLjfa0rIM8xmS26alTw8Z5l8d9AZpfg6LQ+7
Z+Zc7GB7oYXgVW0/wNCwBoGA6SY4PaDBfLyr765aWXYrp0cwFYxGL/D9irR0f0fL
J8/fJFhsT3XUDIAkkn1nBHxqqtoCJ4zwWXTsSbE4uOReghni8Xx9FPIvtmrutfI2
VR7i0Ccu5CoSoT+l2QLR4+Hktu0/h1NtXGSTBZu3K7hhWPPUu7WpoG+fYsWIwDNI
mEOWlYBJCV6Roadwvq8DvwQCzNOQh4qaQBp3sJ5ozS0JSaJe+PKULHBDBS1NvaSH
WDKGxZFRLzGG/f7T6+/Rm7U+otPLHljTLkWaVj9IBWNFC3W7oZkrMirY7Zq6V3Sz
tGzw9oU7eo26YSJKzVrNGL514P2d3NRiaHc6+uePWigV4nGvoIRriiXL/JqqZllv
yGM05UmA7kUF8tgMo2pGLnMfjQt+RzINvtZTSZqDimzUZ6aGFzal8Tpz71xudbDr
F3Lh4X7NB1ijYYVgX6p5T+B+eKwkQzpOt0gLoZywxg2MpuQX5rXAYuBC/ZhWbsL+
+rCeagzIeaVzMRRscrGcXsgN9pTkBhELeaArGxrFowl1jrgBWyIMu6maAaa/oqm1
tsO3hVv7V3g5j3rgCagqU9GyrH+SqRPwjKQjrNX4YXI1bl95fnZ+kcsDmgEvMlQq
5ReLa1eODcHg+HYwYxINAc73oos0AlPlZNMo9VCeh9InA8qvNuWiGsvk7Lh5jk/G
uOeUyrCZyYG9WJDJhG9R/tHnT/aEw+lE8QUTMEV1qEO6kCVwiIWjsNVYlWZOSUdG
+OhYB6slZD/PgDQ8ehfvw9oMpjT+rHAGkKaxzc1515LejhNKmUGvZ7uqrAnJvjgv
sh8N/80angkIKtUEKfOl/LSuVhTK4i7gtm/DJP8vaKtUI+Q3DlwiKnJb45ze/EYZ
s/bqIfsu0Xdfx9fdhmeBL/PHC9MN75Z2qK1WueGVgUL4GkuyzWv/LhBUb8i/m5Pv
fy0Nhyx9HW9c6uRZUONVlhMr6eFmzu9Ed7oBhuDmvsgolPq7k9L0ix+SPNXACiN2
yruFh2GbBL8tyV4+L37TLeCpOumkZEoe4PIw4669xvqO9ub+nvLjPuvHKdNylewx
Jj8PfXfy6UOkcoVrDcmSE7f9w5LrpzI81pRjhEUgHDY3pimVynonkH9QEAoc6ES0
PShvnqWlpHmOJjgzINGQFDYbin+56aLggVSx6C9KgSrFiiVo/bspgnRTpNbapXAx
hDHlAh5KXh5eFNxRgrwNTISOe1f0i53NRQ3PrtHb4yg0vA3wLZ2AQnbbsFqRS8Ss
vpOdPgm80BzK6Z2GA1eeCtZ/8WR5e6xwWfEKAQA8psNYJ2QMjV2aD5GErlE8pNb1
vOLO48O8Z7HVJZe/NM5uwIGueRUWQt3iTY8m7jWzPv7o+29t8GC1T4fLznMLoDGi
F+xxSkGTytf+uB/M0rVbN5d8eot5AFJXVK109dtiZLI+YI9yvGGSBki7MMLvEfZg
GU9qBLT/r7FbYeWOMMoj4XN6wqq+wJspt03wudqryDcH3aEEbeEhRhTCa7Cvk1vL
aT3cpwWuJZRkr1yH6mWuALYKpwasgezhPqJkTFgM8+aoK3qsHQFxuC9/LieTHh3R
Xf5RR9SCv4xhywoVyh0q4NJlQY7GAhAn8nIYoBkdm38hb9SehXv/vLW0sNALD8h2
MBYGK2Ex22E3K7vhAYSf9kquQXhC3dfIjKaHHLgYRjZTZiVrnt6JBlcJbJOCTJO3
KOGPrW9CzszI52Ho/687uq1gJMiL4I1z3Y++3zvhI0uKHERpFmjgbVDV8dEmWIrS
LMKlr/torWUtFZfb8wqL2SjhO0cpX5QKQL/6If9n9flkgQroGyt+PHSHZGPaaYfv
IMahfMT7HqDVhJcrNClfDTXr/gSfv/Lsen8FJM5JCM9qmfEswCcyZqGJtaw5BUaG
QgYj85f1QRShUQHZNDBhJ0rD9uPOfLHgxZ7y9EIHTiqvQr52yOE1QIJmz9hVqLgs
FZkemFdmXNIw8OMGh2hmmP6AQsjMwUIMWil85GsnH+Qjopc3GtttYSkNPm/iASxY
lw4s1gEh3+OKJsSLcr49KAgq7YD8pKjqSFFXcDeAD7I62QztS0JJYutePk8gVcgu
PEvYwgXtGbxMDdBY7LaSy3P+0r6GdZXrbPcF0o74xB//7AfmJxJshWabQAMtjqXf
uJ69jZP6rm3CsJ+bKdUnxbQrjaQRmv+DT+GK80EFyrkgjq3uLS2dsTrLkegctEAW
Wg3TuNKdIvUSjooS3zuhNQLRWYApDnifsHiGJUeGmJR6f/XtPEeF0YutcLbvllsy
i0y8qOaRZF2G9Cz5FT8KagxCeubAqD2WcUUfw8SIFdPVtf9KDK2i+MypquH5SNgT
KHIhTcfhsLa9h1UuBrOYLFL3uhxqUC6u9xGZKi4cfAitRnOQI4ltof49ICAF904X
ZVg8HxS4WWj+rbRRxW5V9FitO5TzKjiXa2/a1XMZtF+obSuT96L1mmooXhGW1lKI
o9hpwbPJLHw5bBuobkH4ygGGaZvhhg++HQyZ+ylZAiMCNnc1XOFdAv9zt/NwUtmc
dHuJnTwZA9obSORw0WjG+x7FXQST5sYbuvufHHZNy5IzC6UUyR+wAQ6QN4DeXMQw
z1ltP/vWXDuu007g/4gDBRfge6cx1eaotgesFWXEUFqfJd3r5Q8zHK9ZhusnLeO+
+URKsi7SwQU1K4GO0uT82F2ZAMyqGV+jAjDnRCeYsKRR6i/YKSfyt0bcFngWRPqY
eKx8SQWtdmGsjLOKV3DnDdtjLw52v/GZkU9byAHM+fLdH2WhuzrT4SePEm1HaslJ
nnkToTrdMaT0S63qzxVXPkgVZ0ciqnrLjNMOSLyfsL0DhzvgI+X+Uz9kr8PaYaBC
VnxAklyxrjiZKpBXcw3aHy25jP7pvycfGv1F+GtF0yDB8S7pbYpSqTtu+E76wCCN
RWE6pklsRTFtWLqKlYHF05AhJS/dhBkgJayXn0yFuX3uEaRoDABiHYSU60Qnjwth
XgIu1D4278bTldRCVGb8TrzfT05CiloaFauf6FbtBLRP7KHuFXgUIULE+7JxJI/0
qnJ/UK7TBgJDzIEHh5Clt3tK4S+LP38m/sjM1zgSkjeuQZ0vYvHd2G1UQAM9a2/6
DzXzFMSuYtZoQ1DeTeOcM2YWYkt+OjdG8fKrh9CqqePKrclHW5cW3zz5nciMt8VH
NYjBswyGHC8VhmMFjnQvppLeXVga8oFVCw7z67kOJIrl+VNPuYBLDqHf8Umm7k6K
0BOIXm6O08aE+fPvNus7gzipgRMk7+75e2KiY2/mSab2sSoCpnJa0WB5ExZvgo4z
XQMfEVTqg4IWik9wOuXiKtLBryzz5EMQgHF8P2DHikUXSUIEirjs5wt/OCLcMPMp
/2T4BTorX6KL7wpivlHlaOIBhyfv+bdWedMtp2YzIe1VtfAIsLRSiSufQFr0ugzT
zh29QZlmkMe0AauseK42kBtXhM6yLChg3bm752pNpLH/RaVnRm2UggcLUsezOJy/
PWEkc/BWdNPkbBTy0OiiRQlCDDuT7b7FpdLVBF9q3DyopA9bYGj9Mmgos54vJf8S
uDK0EJedhgFv6KnqaB3Jco2Y92dNlhfzxRPUQyVPc12tSVpJnIYOWYF3tPIVRdMb
dQrDKVho6RCUKdFIbPDutqjMjVOzjYNYIwCx0fmNUMIYvSn/Ub/C4h5XPq3i5xIT
dc7SK0j10wQxo/gX/FP05amkNAMcNf/je1zxoH4g1+6EwrgWEv9I/dqSdb8IsWz7
+qgfwts0NU0SS95lM69HNcC2SfCbfhKltlHCnAwD02iAHGGiqo77eTg6x4lQYg1W
SdYGG9vYTAMlaHDkpIPZDSHpUcMc8IQiDGOc3aBdbGJN9ZfGFoex/wjg4OnL2yAv
amVBCpSRzEQcYm1gWkjBFlb6DF+OKpaX0W9UV5ilJ7kiMMN3GQK6YLTVxMxy0W58
2Q+eK068k9Yst45vo+p0PId8h7/qUI7PAG8TPf4fB0xoU89tkNfCYZl7N1yqCH6U
5ez6J5X6VvQA4LgXajG5wH/xv5V1dBOCFLeZwIiVazpqguVOIepQP9qmggdf3J2j
riTCixYDJ9aHvys/bFWP36/HzDu2ri51f59mYUSjEKYxNVrF/b7EJUF+PX7atyTp
bovxxSkgLf3H8kJIIhHpBiaKThnLdxxRujtNj/+kZAOERQHpAVN3w9poHqciIgtY
YkGMtWPKsRXNBI/IolX+59GuQKjBcQej0Ggv7x+iQXT0w8VxPcYmhO7rGt3p+aPx
AfGynF0ckwI5SZIBG3eqPQdhsRX82Q7NIiN7Va55l5fKumzySQPGBbAu1Vgcg2/r
ipZGxPWyGwJ1cmFhNyF4o2IgyFUEt7ZPEP+7gv5lwIWxskN2Bfvdm28FKCCCqtoh
bY3bL4P2hq6ZqdNUQyVzR8me1NBWvd2AMNuEUDg1odaMmVFOgwTLPxK0KrnbVs/V
wmfPStvLRo0IeTHk90t1w09gu0MFQ4b+cr3vkgJoHeNAEZOIro+RbgjCsHqWDQYy
Ikp1wcnPyRa6J1/+qzmrq1nUtWjIRp/kEabwIY3NTMK7ajKV24wcVldOiTbEL7bv
ZVse3hkja4KOCX1iCIGuQr+jFQokt3sWLaosKPdeBV5MWEr+d1E5mzf+0uAmQTEH
BjkxlXoKVNhqrw3WZUxs/9ZRMHVVrvoMudGzlMdKPkPc9nGBLbhU1z3WVGUnQWHj
Bw6O64vXa82Y9nHsKXPUMAfZamKepBdLjUUHmznpjGC88ciGmSndPv7DYKUkWwZe
pOz9Rj4BTemK3Z1dZ4+Ffl6YPos1MFTbrZwZpvz0cMYMux0ncYbXV6mAcImeRrgb
qtH5oQDMwUN9iR0qyOq8EUg38DnAOJYTKiVPNU9ZqwNofRgniE8UnSrQQF49gf4W
dzgX8Uq1WMNFxU7ijGFqK76cZXfo93w9sjCczVaPtN4XjMyQWDiqBiMdTLE876g5
/KYmjEd6eJOaxUyJ3iwaDiPpjYBQdZILxCJC3OlRWOvr1egoS2dEcOVUlw68h6ez
HLjHsBAj7svwTu5BpJluO12RnLzLeUETItQd3rldw3oW8gljIpfQ3WYYvdCawGqw
sO6/xjPu86Aj9+VgXR1qLNyup4zWawOWJ9easXPUjxWIXcjntIYV1k7xZf2myYJ2
H286HBpUwu5V7CzmbFrEtzsN0yblDHi3XM7Tkemg8gfzIAg4it8dur9YVciYuCLt
iUEHfTZUiJe57mSzafsCr5+NucDXhfDlKqYvpqqYbizVWwbrq9+GVyJBWEGYSkzr
gF5qf0h4ngv3TDUkckOXUreJiToJ1/RwV3VLM9yiMg96WKDile8dzW65Ze8JJENh
O6G0dTSVurBZSPHjxGKTOQB+xtikLVZLpqpGaeiVxR2OMr6KnrqRi/WekFnT4Ump
jePegGy0lN15Xz7Yxwpf29Li/an0Y47gJ6kXzwma/H8I6sFyt1XfozXBV5ZY3EFw
UPbHf99VQMv+RI+fujNvZnTINTCe7EbLKBlAX/GQ02R/E6Dgo06VXGiUtJvWQd/G
5Zg6rQEjpY1SnSlfhsJrPfTkbQp66qjyFFZuBS1kWhKi20xSlfzy3BSjrL6bbAom
vFKVBs9yBhFj55+2g6mmwaQWXa2T/MZ+/A4Bgj7NrIcg8cfpDh7NtAwPOddmu9Q5
V3Vf+i5siSaljnABsb5SHvOFaAcYTBxFXDqrJ4UaWfrDaeMRtaogi8FnxMstdAPp
mODeRs/jm3/CvJyGI1Rc7TnE9bCdD7Bdx5nACeyfbgVrJYsSvsU73ZcDMcnFvH0r
X1G32YKgLvdykHCA/Nw2sN+mJymEMoIthLMUXkFR7hmhRi00orYgwvJgZL0ATEY6
H6cqNOD754wZZ1paePQX8bNWB+2WIs4NN6LWul1sMAdztfL4U27kEDlwByy06OXC
77ci2MI1K+BG3JilnyZ2mavQK5LdNziEweeSHuyKqAwYkaBqWN9twHUT+7FXPr9v
iiiUZh4/h4leQiPiMxYJIyiLAq+a4O2CB33TIliKV5p+5YEqae0EaqbaxodsAV2P
FOor5IINv0LdhxXo5mTn/nvp7CriRHaz8F37DM/fZx9t6kJhahWOCf+Br/6FoRXY
63FhxCe8KZ4601CKGM946uFpHfjpLK9AqiRxLK85tNGCrGdkPK2urK6xZf9YUZOB
QC3FmLG8w0L0J+cHlHLS7OKB+E1PDFP4vpGr8ly/K4fKIcnKEJX+q/pxS38H8Iq6
w1VCGOl1X7RJ87IX+4XCN/ptzoP6Q6Z4rVhoi5ce3LqhQrd8Qrwd+ODOiNH9aEia
AwkLSu1ASUB/bNSUSK34sLLPfQcBiCUudz0e9UKIoUKv3bgk9ydIJrCLiFX/LD2t
MT7UlygVHq/hkNyBkxLtr3fG+YMvwuGpl+mJiKFT8U53ZJ71wWmaPQM4a/D24zai
WglIkyTDGAe+357/ni1IpiJ8p22PPLq32r/1+ebVU9Fg5BQhlXjbqJY5H5cf/bvK
KfdlaSZ8dXYnZpuq9FIcCmvUddl0kS065/S1wQbJ9yTE9j81il0gj7P2OQKe4Myr
JfFI/EGvhXfRhDaEqufyBZ5vPwt0fbDqqRtLYxBIM+C3zUwjp+v2BI77e3XGBMC2
4ACa+qLNpjOGdAk7KWErj2TPiINAiWSTliFoW6J/nSIduyaS1u5hN1oO5trG3MGJ
h4ds1xKbxnEexFKx/tx92Ub6KZAkuVWIE/r9B1hyKOOBt48mVJPdwzYNHTOIHl8Z
mD5NEOlu9wRf6DL/c2SF917lwWhmAxzbw/vQJ4FnzP2u2RE2NjyWnWGuan5vCnw+
sJTB9MlCRLNnsQ+eTkQy2syMxvzyG44NvomwB9rWZ9PV+t2nysdT3UyOfhylpNaB
nAhZhnAHwYhv/2W/rjJoaLZqvEADfyRuI/Ai8+enG6toaz6Ot8iJ9bbUyiUlnD6Q
mIYrjos5YdcuNPL5owHw5m2Dw0/tS+CIk/QMVUzlg79S1pflJ4lxLgE5RaPitly6
Twr1D6d1YdZErpId6TpGtuwTJgTihwfp6wmNm9DN9BMSeY42zhOLwlN2cdTo5iYG
nw/tyEaCqpNSaanvrwXN6h7bXLrOaJIhua6DmfO5BLJifLYED7sRoLBf77jODfb4
C+SLJux4PH8zvUc0Sq5s5GfbO3iGdcN1aMwn/j+9fzf20ugZzaLd/yNE9UcHAjQi
f9lSJyEeI7WjdeFHZ+suLkvUVxulnCeMCI3ID0Lqym0ZU/dRJWw4zq8drmXLILYE
sNOarYqaCSiTTzrb0OZQy3CE6QzmYyFIg/lCwwM6ZBYEqcf5ijLCQ6f4IVp36sfN
L3YtaWA0fb4Ck3k9LTglT8mfBWa6jxG4YRnQo0MXQqXNRO1SY1aHWxVcoZaxctPl
ouEFztmWkETuArziiWgKQeF1jKJ06xflmJdM8UWcPJ5+RdSDdBCcXHlNXQXQREgf
I6IybhlDkmGgaMLfq+w2vylMXbQgvRK0/QhNIjRLzSDBQwxhAPAdUoWaEVcCforx
2gKfL8uRRtiXFpOXROGlLR59cmdNQ7SqaSsgcbkvfd9nl5nF6dpf7hfzqUgTg6Lx
tFRWZzGpujBBPyjE22VEbyehZgFuCzxqUTA22OtshPoSylFx7ooRYnUlWxk3ViSq
Pm6vsCRh6rKgD4xYD9TvarGdNWHDO6qVOLxOwVdh+91D4zuUQNAYCpCT4bDYXFmY
KlKznlKr1ce9E+g8gdVUzJgECIN959rGzmiQ5R0AP+QVu5VxGStNFYlujdK/ZKKG
6EsS9wIwteGM+BJ4/tQWWVOTpTBx6AIxqAlLJRlXBT65JzHcBbymTbAhxRCrs8cd
2oe7x3FQUrJnl1O5H/UVUkti3b2f9SXcXLs46kBhmpv/J0+Cm9LjaopJ3/+zHAX9
PzdTj/B6uSmacVxYxfvuCKkadT+67e8yj3Uyj6wgpTUgBCQLxErhF+wDTqFTxgIr
1DUUmD85d5E/bC3KpqoAQkjI51pJDyVCO7OymETi0f481zhuTL/toOUALNQ3E7Mi
M9dqAMPh3lyflPslrRA7QVI7o4B83Xx2817w1+Bpndgzpjq3yPou/9nLe8cCSEpZ
OYwSnWCkYntIWMNHhtP9iLCUIJQs5Z7v9+OJC3ytA7U507RWMICR0fEviu/Ko9aC
gA7qDpE75Q0QAUyamkJ6WNyIiYUNNqD0ociWZbH4tAmwF955sswSZmMjoKVkCy8P
W+eYjLtdZ8gbyN01DWqxepj9uoMwkt7kaGT9SQWtr6QweVJQIKmsLdzI7161A3wG
eZiN1wYgj2i9Q73v/CJht+v0zRfdBXAO/Kynz+ItBMOQk73EqpP8Myabf2zL/ueC
swEh0pFn0/ZPhH0ruPrHl6NLiZaQbOIF0xyC0TbFBlBNXyiUYSf8zmOCx9dNbU77
rj+LxHVsr+kGb43eBpNaHlM41+W8L+DBIngMF5Ts0Qjm+GTq2G1DVFY2eKTWB29V
ZA/1hP8j2q3fUare6UXM3o9jQJQ9mwbaS3kxyEpPCycRI4UmBPzotCMJluTWi7lu
zsTEe0JHhmXwPWcart6lHmTS47K02Jly04sZZ4GnbcnupQHWwXF1D3lLg1ej2FlG
sQu8b82kV2dr6vIDRuwc+mTqoEwaVJKawRYMzryGRYVZQaceENYtDnAy04k1Momz
SxSIrQuvhfII9C26u2C2GvdSyop47Sn/4BgBLRw/I6xgnEHS+y6bNo76ofSnzBQ3
+7yKClOxsvXiQNNHdrOY9TO/BVXPhrpQ1S24Tyaw+dr4LYEmI6ibE5W27lRFXoTu
gMbwR97WGEEWdDVRsv3nHPbgiMtcMTk60JPeiNxZS4XGnyAzKr/FMXftGr6cq9zg
V6C1aph+bHlhExcRodLPLxUc8JQ+ODW2Y0HExoM9fer2YPxnNee+lhAFNU84fA6a
dkMWD5XfLVh6NtfoZOLXTVdHCUfhAg9VJQh9s90klFkQT+J+W0h0/Xnl8fhSOGSE
orffaKKA8lqFPhsuGSxvSehKgX7kqDOaT1ApPGhg77gBXg9pA+RB4XL/3Oh03v05
jRO7QnlkJfWqPA9cgflscv9P3d/Qu/ZWxklhpCbp4jo755ceDNCGAcVruZxV2671
fIQDK/ZgVXTSJ0EBzfU6d9Jbm/39vWi2OMkMkB7yhcc6XaLjcVXCfCmgZFDINqcl
aaPOs1DcYvp0Cs9o+uIu9sLT3+boDb49Y8gzngp+ogTsQ7NXkKGVSc3d3RSKJW+2
Lcj9a3d/G5tqf4z4pcpxmj1WO0SYJ47KcU6nhi160shB98u0HeonpSiYA4zXDRlW
w539HXeWp0HsVD3X6sMUgrz2L7zelVEh1q1WlspAY+OITpViHi8lGiZ1XC4yviCq
ym9D6PQRde6cLYeJ+8jKWcnR6lUvbNgC7ya5T+PDLFJMe8hX4BIQsFGSGVjs4eZd
uuPkc12VmF0kw/4FOx2QZiLg+bSECTDFiDWdn2ShoMFohaNn3+gg2XQl3hDrTUx+
N3t1mPCwAIrex6daGo7IIcH0H+qxUq1/S+EaR9xnH1Q0UrUlEbaJsGuBJgl0sFvu
cuZoR09XfHA2MhYj+Ct0bvW58SfO7zdt6AsweMubbJnf/82LNOSw9pOTNeknKUGN
d7jL544Tm0QB+C2r9LSTUKWhQd8HdoTxVEUUOa6mQxPAweyavbFLn44oVb+7u18g
fshyCfWKXPT0I0eUBoZQW8le3aM1c9BHxzkKMA4pxxAphjJNi3+mjmBo6sniMPSF
euFaAdsPVmW8UUw/fuyya0M19iylizCodFWCd35PLy7gRFjQ53NQWgr62cP27rwm
ixKilFNHzHbhqorEwwgicMracdomtcuUvPxFt11b4jhYuZp/3dGC+nFCGCVoXoye
t9PkfvzPHfeo3b7ao29N5vMyJAiZ/mwaw9cLoaBh+hfpTB6V2ZswK3WCoCJ1bJi1
kKECZj6DgpnTK0cO6MTfrC61tFoEkv2fmczYS20WUjPRwcSwSV611ejLnxgFlHgk
CI8H/iL3J6YnVyqeLRA1sQ1nNWog6NpE7iCxNinYy6Umht2wQpLA7sA9SR52V5Hw
JzBoKlMQPEO4XIYNLdorhA788dd8EFVtax78c/i3km0CRFmVizsOe0kgNH3VgSrQ
y+kU6fxC0qEP0bZJ0RSHMpGRtNPu5mz5/4pk3VcCbrvW2KviGlX0/HP6lP+RCLPk
+xImdYljvrWnIOJwSOdakOZG056ZpNWe4Hlx104XgxGPSWDKK2MIrluSBa9zyCH9
5D9SvMhSGUsUZy/c0xZmE4+8U1SBgh8sMhsXnbzoSPK0IvwGWXUJRIEHOWjDDBIz
iTP5UfamEQUyZMjFSOxc1BqyXTbC7/Utls0oP8lWpZ+07X8mDiofupSPrnmx6ts7
vkERiHshX1QxHpnhSSiwzZTkpaDH7g6emIxV1sf2ACqMxXMyUHZpK6FUAOeDVFMk
4ul2PdS5J0z5LgcKzNt4T7xW/IcsO5hccuT8HKKqWqDqOJO3P/UsdS0uYIh1Y4HG
JbgH+gm9uy8OY99qKveRBNupyYaxdnvm22iC7DoD3wjmpnyDpV5EQZcM/KWODt1j
EmHkZeuJQ2ZzpEU/IgZnKhMg0Scjf6lqg40LFE7Jd+uIpiFLAUnJzS6y5zFxjDoY
buGzvcHZf8v9JnzdjnOHQg4SI7MO9FOc3N1Va649INEC509DM+w0V5tRJbvCWfvE
b8kkHf0EYrLduyWvvf1JqnGBD/Fw51XkyA/6m6kKxaPc/ONI/rXjS+I0odUmq0dd
IPPtJlqzdSaO90a7w+xLhw1JsHRpLe7cQ7tUkWGxBUdGweUSJfb2ikXgz3HEw96m
OW1Gv7gCcXtwgu2dobWsCIN4TRzza19Mk1CbRL6EZRB+vg/em6SWwFubPTBN961j
cNgfyz0ce1Q/M/9TmQ2P8PK5k5kaHDR/f4o9Z4X8BJEwQ6yKWzLkxPrpLSDjzveZ
RDTCcDCtyHcrBxOv9T9P+AH++flSd+ULN4ZoAwd3OePum/dXNLozoSjyo0dTiPIa
40Fwro35F6L9XGAdT5diY78TGzvprMTU7kVrXwrkVEjjKOKlLSTy+RD/GXm+6xaz
5K0Nya5QfwAPXtoeu7w7stVmPA4K0hn3qDRCnJvFf2QdiiBca/k340LMIP6usKUp
AumYkvsQnRHrnJdd6lathyknUijNjNKtLvh0WS/84K4uobLZm+CKaYxFJ5En+cfN
ehNEv8pThgx0DHe81k175rCqQ7FnuVo2TrzDQt41wqgUwvOJf2Fvl3ALzYRyECZ6
uNpzEHQxutGyDv0g9LW8kVPEg3ptmcCvq7q/ZocQuO7CN5OScdLrZaJYd72Oy+OA
w2lUXXGqm88327cPQeA8B6Nz0hosWTXTppbovG8JEhXCBh9zWEBrwj4/JZxRE3+C
`pragma protect end_protected
