// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:38:01 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
J7muSFWy+CDR3oVlOcXZzPV9sIBpCnr0xSS6M0Raxoik6tcFjp072uv0zxtDE+OA
x+1l09n09NCoe0ZoZ0Lv5H30o3ePQ6e4HOM2YEvSBYBdHS5lxiJPxJ6ryXDh5wDl
OK4apiEnC9T+ARgYa0Wmbb7c/kjcvcDtJrnBEItML48=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8352)
KfnOJSMHEEheKyQqqzKnZJFLkopUeUFARJ+GxsCsrCQoxYbOSTjUgNXd9KpvUc6O
iV+7JPhb+z22hT9tpBtCE7qSXN0fhw4ZXx1hNZ+EIxqjZUOPb0qbVTeSO+z5Vp3R
HVyyEfKEBvm3V1w8RVU+cBRZJv4wMJyOLLaVxkwLIJa8IB2AWeSmyTR2TWPgI4wj
RIaN5txeSiG684HP4sHeSw7JMi15u6Lvb6AHGfdOdGzHjz0PLxQNHAjmH2FoJaVi
MilTvFnleDvwLdTQeK0ntCHzSU/ZZZtTJ1CMsJyh9M7ApK48aXpktPYKC9WYKHU1
wJaHnKHxoV7I4ajA7gAFRjClDWkIauE1NsNa5ePFVpSetkEoK888GxsWs0diTN/T
AJkzWT2JB6cKTi2PzNAIQByRNfkKtvPBGKpkKVgYTqmK6NmhA+AZGKBztmrPAS6d
7iy9GFooLHHFYDUEqW0bLL+/Yhr7f1ZdYvr5I3Ph79bXlkdKfQxIPz9i7chTiO5q
2YBy43uT021aW2U7vkvVhUgdqq9T//lzBzVDtMt76GMjfsezkBo+0C0OWAAIbpqO
0bAbU04JZTBW3lwoFlYZQmFIKp1MXub+aURqyUveu1rQsp4RlEvEceNHIUD9dT5S
ULAGi+dAoGubl2W0NFeouNvtA2yH8P00YhRWr6LAobO6k7qbInCHnt4hUMcSHO0/
WpVPfgUKO82GdrIKrpu3ZmLfVFvZ3HoejFVG8Bn7x+mCWMDE0HCgCypvRJ0jR+pj
uJKKKUH9bKvLvtWQdmUaK9BOg/H4bSNDI75o8YNtCGt+f3QmgoElUZZi7oHeXTvy
jhZti0qf71Wy90v3vebgJDjoGBjOXpGdoQKrozThxuojG7wEidOtrejRNgVD7Yvu
dfbKo1oMoEgN/S2EEtebDwRr1AvfuOpEcfAXlVxmw5MirdQtVHKoNvgwEbglsLyj
NILIRCn7PmVVZDLue5y5vRepW7/a/UqO0S8GgjZkr/m/t5J+le4N9QthuxH06nUB
3/VzJqnkIv3Q+HxzWkOYYqEFH11DnyzFbCMsTsHGf/lfuaiHvTpQovOP7a8wheiz
/n6oZk98dMlXpNVtJl6PWJ3WGJPKwYisGOnaJoq3AStyCYwE3Pet6lA94gt5Sza8
+633UetEVACQOuhu4aNn2GfElWQibCpDhbByuaj4ibMFC4dUXcJA7JgJifiCqxD0
k2+61Ry5CaOSukdDy8fBUFzb789mn5yOcKDOyedVsQ5bW9ud/D1QGZK9MnaDBQLv
4utLO89xJ0qdyCP1jlCkjR1iBmOgMqvNuDbCDpz3TVYFSshcHYuAB41/R29R69ZC
8nby86jSGqMpShYUicJGzSesxcJqSSLAypCADWIZj792d20t89VGXMvnQkkrVz/z
DFrrEZWOr7bZ5pXnGLPUMun8LmQY3hnSzsi4lS9UAVC9Br2spIy8+zRb83Enq5YI
k23IO6tAcmQ0fwJxf1rSWgghY6T2f3oS9LfEPXVc1vfjEEZR175qvLJ2PIKspnIL
9nfuzBCt/CtNHU1A124QSLDuHLAv4h/zb7ABLHF+8AkhWzQ9cXg5EhqOy8RSPpL2
pIjPdiAheV6LOTp6Lmtoa18fl/GUnoY9hBR7g5Yj/piM0ieFgX8Zc1OuOFKtLJ3e
45pSXYNbKHdiDEPhMR5qoSG3VPugdkhg88EI376VE482N5dQCPUjZ9yXaY8bZQuk
eysk2+n9fns6Zti122F2T0lwZR+3tsinAEN8hl843Wg8BKrqx3kLhSCirLKPGo4C
Yzqb19VSz62XGukwF01cLYu1AV+PeR4dcI2iaguYk3b9J3a6PKfTN/f0tQt9uTC0
xRyvigGzBqcdQq51GR55ncmJdKfFKeMy7JOVjHpkE+3rjnVuEHrQvjTHYmtVPZoA
mt60Ob33YCz/w9WuRwf/5QHqSxgTbd3gwzmHs5bVNJhD32yh7jrd/vpq7NapZu54
B8hQ+DIY0XEVxrJofxH3xElC8p3v1A4un/4QYg9ahqX2JrD7xYU3aFidl2OdVXF7
nvvAkMlKixbQnFuzr4Ff65COYMhZRwcOJwz3MkPLMWt3OWi/ksgFe8Q3fjOl8NGk
Nkn6nxfePnewRTzd6eQbSX+cm1WVDYMo3ThJ5aC1nLSMPcEw6WOxTbaPqvbR4GyN
zx+WE7WJV63/45F8ZS6qn54jRQSWiM9nlwBugZND5TXqX9CyZkYQ6aLOzir0qi4A
O0h9c4xqN0V0z3NMl4A0eAVsjA+m/9UGPVJeTpAhMQDlaLvaVRek2OFjJd+nkPX3
7gosSwiuxWQ/vH1EpRpIOFVv4+KwN5EqmVe1fMzBqZKYpo6tir0sDVgBYQyjY5y3
oRcDDIkkKv0KirtpKw8x4NSYU0wJfft6Xyy2x30XJnO4mPZVsILF9fhd6HwE3Y0D
DjwqTWPiRoaCSGzWAbEd8yqN15bGOUUVuxiZ0Kf0CXG1+WCnE1mdu0SLY4ggPfmp
jWGzl1GiZ3Vm2uAyYCFfggOhD6AsyU6CP0OaT33g3Y47ZOIzlXCCUCb90MVZ3x4E
Ua/zfWQP1fsYVG9JHeWb3hREm+RDDVypRhswPGI/37Dm4s9rvvB2Z9o/5hfkxkuA
syD4vOjgEx+wAXcuJ49dRSjLWZp1Dwe9/wjmQd+wwBxeTLTFu4/b9aCiHDa6/QSN
qnA0+Q/LtM6hCQu5K4Ovo8kLvreo9c8N9HBT2PT7IDDbtOxHvYL9Y96ysOwgw2nZ
a/V5rS9yVXnt6GvSxdoiSfgGfgvjurR+XYPvv5UQlksWP6AdYv8OFOXH98TeMmEM
NFSwoRkHW7an7+tQrDyKkvikZf8NduHpUmkdhHXgeHynTtN/Jtga2VxnieZWVj17
qQ2Uf9820lfjeoOjv0BEJmshOl08G+DSQ84g+YPw4PjSHIcOo5MVL3JF+AUk8ksN
PIvlH7JS/h7SqZTsCzVDURt8LY0jnpPq9kr25WX4tsz6l84Kcyp0zQs48g0GRr3r
+AYdJR73pNscykKttsAMW/WpsaMUbcl/G3TrzDPA0tngJ3AOHW2K6jcW0nbhDN5r
KZiyF8dyw2vLzhexMgtQhviNNmL85ZPr3nj62z0quxoKKIzVWSpJGze9UXlqmMsz
ajyeTTHI6p6sILr0n5fCPuYGep4RtvQH0iW7D2GJa0WiYz9biACyfu4PxdzPOD3x
m+4dt81RwBmDb9aBni0m3tXETZpa98o4aIY7WfiD0Jl5q0z/AJ38cS+75zlIkih5
Qf/JOSeQ8YVqno6HGbM/ckaua/gr9FCAz8garP2hkx7oWHZdTcYOFMHg55AUdHUH
6rixAT/c+HBxEtr1HIZ3jmkOlV7FFBZdWtS7NlsBN3CC8WFiK9q7NoFRMOyFWEHN
cmT62OYHxCd/n2mnKFD1JovHJLSNQ5hvVyr0owvgiRLPjXCYFkToGU4uHAAQF1d1
h6YFMDDgwMp4DThZX9C98Zkfku1T3+hQNamqMwfR3xW2rVAtiDJUOS7Eh2jXjLLb
mvvHgE/QkczIJ6IOg2b5/SJLX2pkaXrN3tWCMr5PwMDdQ2RDM22zBBeKBrCa8YaL
2QVPuwzeRvXNkk+FyQ7Vx/GjaSuRQUaQ8NorVNrDq9CCaMXFOT8zml65IArcej52
mMhuj9Shu0SgD2GSs0+7Mb1GZvtDUBU2oCUb/LQQx/kCBWrHHVLddRcVGnfPGJdm
xARx4M88Ne77jc+yFBrCM8zY953N+mz4oYH3QzOlexfgWs5CDQlD3dWNoC0coql+
mhZFx8qL8OvYFwKbKL3a1hhar4N8xLXneTsY3DNdVn2M6xV/1mJKaNuO6ECNL5o1
hXy5a/wsm39ovU4etUWRjSauB3mMKDu3mJnQEE27Kk3m1VSwGX8OmQM2eb3AouBv
I35NdZ3z9dfrLxCjKTTbgR/lI4mUhSwQn0Mw5EOHUX5YS7KhtZCQXZfZBUzN8xv1
qFFUzlqfNpXgHe29vKiwLI/jkxJvdrjFcL3D2Qn+bCaJ6m1iEf7xu3IV84FiC4ia
imly9UzVjAEwOfn8sEYqoJLpPvdZnJm1uBxQVDOa7kKt7PtIpVR+gh+ZwMFE5lYP
auulYYCp1gwRmpSlnzktyNVau3HcqF58gzy9tt42FuvkquElyCcGTh1K6JbFxubf
jhfo75dpEeitEXlLFhYY24YdH9inYfIcqnCzq7W7OsMtRbUb2IahOQjnZp0DO9jF
zjB3bycgOYY9Ch/zXQu2OJZEtxmQb8rhgoP6ECHlOgaWy7tHXYZf6CLN9IHCrz9a
YVbGrDEmW7NNzEdAPexE7DOIktVx9zoEEHzBtOLAclXvmt7GJeD7CC296ntVbBr4
hDiAtx5YFoM4gqrgCWDnAX6/OZT9rpouJqvSSKeu8Uxd1GiFJLSVhEjL4gFSnL90
HiIzNHm9Na0EAdchsetL2wlHObs37YM9wcZ3Xt2erR0f+mVeGxxM6uYKqTBo0Usp
/L99cCOjdYxcsFjF9hsO+5wLSKgfit56ZuePJxJXF6XmY7nJBj16Xd6dH0l8T2cO
56Fymm4gRuAtHtmEYMBGbSrNjfZDYb9Rolh0FslugzQ+arvELZyeOE2Hg6nhha6Q
YAANrOaXqMiUab2i82/v2YFWdvSy983m44tIjJ9aU4OqaEBOtlcQmidnVRyy7jqB
WdDXFZjEezWjNWgHZ95l6WJCeBUi9B/gu88cNoZthgSMtcA5WZkN9QaqC5Vx3hHX
6cSsYDVSHY0AalTESj8fFOlOWt+nLBOQs+KWhC/lKxbdJ+s+WL9Krbsq3T8e3awl
1GOtJaQNm9PshCEBqWrujzJ/bVEefRvhuy2vrjDqRH9j8j/cMESMOW5dA+zrMmhb
zgyTEeVcmAXKk42cq9ZlRXkoMjHAzQMXhvVoWlcd396q3sgtiryaLy6lQnU1KUkK
LrKzXYHGp0L+Wlqhb3Nh2F6jHU14aBomqCEH+GAiXo12BCXmTHxtPIwc4J9ENMds
TzLQPK5onQNwqSFuty3NsMcn2ijLcpsxtg9SB9PNMBe/E1opdbCDBjVB/9GGysN+
7m+YyuGXmw94H78Ya8XTPsQXu/zJNCgYMS5Y4v7Dabx/+MJiI+xrpU0IrpjjCZ2D
nn5wcLx0f2YDf28a2oeY+nhEd2LSuOzwcH9Ew/HBwyamdAoDmYJKVCLcZpqIdaWG
2rx9mPD4aE/S66hElzTfv695URUuRuXwBf7lnk4wvkAtUSrjt6ZBr/K06R+eGYfx
Dp4lB06moRMrVSRdN4O5iJGPls9EImGqs+DlO1yAeWXzxtWtakNBooeC0xuTOlXq
zjfZNTtoq1xvZ+NF+EnEZAkTQ6YB92IaeQZbbNZFgPSI0mLaIgY0RjBM/+dkdFun
E+LCPDQHlxn9tGZ7GQxZLGIgmqUJdeWST1+IXTGUpVnejoNXU6fJACUM1+WGtnzy
pG32Wu+vW3plLhzvpvxZ1hC1xTsulUbwoyyozfNlrj1pYVNZgGBxqp6o+k6e1lEz
/NhTJjgxwn9u3+DR5vYGxmde0jGiSK9TBYBcIVjDQx02wqy2SbcdXgEDbymXBcEF
7WT1LE+kuJgvBWuoM7XA7G/G2MiRyP5ux9bftO0ikjBlrM6mQtXuPFGtBiLdlxhz
bE6c6ZVHxCYf5ssoId7x9c4Gh1nV7GhGK01DWZaqKU0RQdqm7Zxg2/+AuPhPAvQb
ZFgMSlczu+5MpP+Q5qfWczlrxkhbkz27COs6TO2nITJPIuZ/XoYH0qWVB/g87/dv
DLq5CbCoRX2k4hk5J9Tyb91EVhadHDGVkS6CC3d4w+lUwP1ktMY1DGlLX3zgtAzU
Hodye6DyL+HTwDQN7wGXOa03/1z/ONkHT0KG2zaANyGvso0Zd7odtFrt/jdc2nLd
lw4Nqx9/EPxgPiQKL4qg9Ikhtp2Nc6WM/fglEfoNXB6XRVDvuOqxHx9tljJoai4c
muF9i8MON5IKPc3UeIs/9qqXIBMPyjuGZBickeWhaDmn9I8ABOMUYv1UybeaGmaA
XK/+5e4GRY0+GyurtYDns8keN2hK6/ZwKxzHfzTcNDFUvCN368hvdAytzrqnT905
Mb+xPff4L7B+xOWt7o3QlG2B2W4hP3S0HY4m5tBKm99lOsYgasKgcc/K/fwx0ib0
GS0K3cs8DxK4ZUapGCrcuN2WGNmFGm0i8NAIZ3VOz1UbyHrRBzg0XzJT4JJM/PoA
K5NF/GvyMe8QgHt6k2NiLQyAbtNHFQdbT0nAP2YVcYx6Vu6EYuN8NV5iiEf+O5M/
hOobzVa5YSKQfXqvYZPwbMNIKnkeqycBtDHoCzltzEN8TYU243oRYi6sldlLshae
xvPjayKQmzxwaDz5fp/znebvSwwzedDL+FhEDKOd96iTJg76qFi92yRvKCCzPb1X
C5jpSypc05QBwo9ALW5D14dR3lSnGaWA/6Tx4lWVyiTvbSYBuk39cV5p/YSiE8Ya
fxaEkjqnWG64x+F/bOINNQuhq94DmS7MeecEH8xGHSC9vNxB/CsI3koZnpT2azEX
8uba4LgfxBzJfM/hG4d6ygdgAPluVVZdv3kYTb30DD79zs3b7b0fURSjRWnYS4cL
6BQ7495qid4Dlyd1yWFlkOvU9aJIilVi019hqO73bEDy916k4Afd8hePhWSuKIpw
C6iamsBYDOgPKTiZEywZZTOywp67JIycCC/cODKRy9MnA+zGbdtUgY8bchrUW6Yv
VVxucvOtj3Hi8JdVm/aBTV4MD8dC6a5dEnksE9OFKkJ7/E/OB2tukOmdUZAkd4NT
z90L8ASyhrKUK/gi5TqeyUHeCGshGt9BfoSR3mSDPFb7oyL5T2xek7dCamal2JfS
yxyTmhT8/jwzAkv96TVEjlZ127mKe9dygDZxlOam56uO23qr3+Hzk+hDBvg/8eaH
AXG1NEJDr1bXZ+Lvoqop/zNoLBT9F91+1fCfa0/Q/elEN/M0E3nmea/lrolq9PwT
V38//raM3Aeq7ghYQQgfVaPC1X0h0uPKkv2/BwlpPu9r6XOlT44MqQWMjy4vvI6A
xg5KkW2imR7du/W7XVHyenMwOHf5cOAa6KKnODB9PBQ8qdkh5BKlgTirKZ/eMCc+
cQMicoRRn208zyGHpxkCM7CLjXImmlmc9/WqGiyadFkql9rVLUuT9NTx2zvw7Dxb
SVNvqwCSqg7c2dZ9e4lBSK/1STjbJZE0Riq5gn3sbBNOfmr1PftsJvFO29Ma4y0w
peRkbZ4Imx5dr5fn/pESzJtCmYz+oCL123vYHAPOAj+hF6ZzG/7C4vY84cJJcTmy
QssxudsF5nTV7SfoVu2JA7/HXJ04w+X3BEJo8LbKhOAoGqmTYelrZhjoYtQ3AB7V
hpni6GcVsJRZCtnTf+EMi6RU5cSh5JVAhLesUawmt+LAF2Ev7Y92JI22ctoE/eu8
fXcSKAAkrY2KXtbLmIJda0oF9dlWZnli0OKZ6vqpZvl9S3uobdOe+ZELLGGR8TBr
zbtI+7fx47aQbdtt1/7vU13n1m1OgHNjE4H4Ci3KWawE2fZzb3gmawr0MeEmAZIt
S36TR+xd7Tu5JNMQ5/5UHzQ1+aFBtn4GJN+mRtNjvwM86SPL2+Qz7dBVR67g1bjI
xkcit80SDGxdZl0vop3NIc28rMS90et3EnAUxuLpdNN1IqWi8e0DuNwiZpuU2PDP
VykiCFP3Cmy1d+B9xpoQwTHzR7qfA1vfwmaEd1mLD6HkdvGQpvWKdRfF4tZfaikK
p+Gx5/j0rUIJAX0XmbN6z6IYI78KbSXYBcD6SpajdrviVYOzdjTYIUpKXw6vk2dw
k2vkcgpqeiB6XfrYY96OxWlrA91gvVOvi0En6RSMllPNdGQM4d9TC6T8DZT6ZHGM
4YizKe2Ok8mRVDBMV8S2/AxEqg5QeQMWusZbdQhW6qqmxNscOKIf8SWDJp0s1dqh
hiDr3RyNrnOh12bu8LzMwijeHhb0yi0ZofkrNFl7R6RisTERIBBZzG5ZxLZOPXBv
jNkjPICsbiWuQ9R/v0u27rXfl0b6Pm/si4HgItYCCwJvXwqOauoTjeAnXNM9XnVd
SG1aL49c9uvJD2dDEaq+inodo2BbN+TcKBXxF5AvEMFCqsniLsFBUe+a4xw5FPlm
gy63W2VpBd4hLHzEtYXOy01CqSM577EIPug0pEzrhRBzeZ+SPETuAc9O5UkFfe+G
kXB5bNEOsJUFw7l1MCYIHAjGkOwM1XstIH/vN0lQ+yo6JY08zgfEdEO2hMdKu+va
fW0iovHqedjp+47W3SdRAbsWJKLdln6k3tReBaH3arXTfvJTowgMWah2O3T98uvh
1yRZuEg/VH4W794pinQ1EwEXJmTvUAiMLZ8RrauRB+WmtpB52D/HARQxR+Q9qwHR
kyn9ncKQsAblA1El2/aHOeSTSRLssSy7UM7W8h/0kO7CpXERUovDwTySOPonU1JK
iO0cHOmBivuHL6mzbvsElMkI1B9by2k8hwrZHgdxZRARcX0OmOHGpzrhSdNYJWtd
SyL4YN6w5IQ4CN8ttEwvIEPWWRw4q/JaFlebWh5j50mua2IyaoozEkinVbinZqrf
6XlHesSjTNj6Hzsju14BO3l6bO7aQfZ8Zmkkq70J+z0gVSiNYh7w+taTm+rhT9iW
1wApHZVgBxD6deB+uPq1zJQp6KCNygTG6ZpoP1VOWzv+/il0L0j7Nb5AmwLDi1+h
2bwgYvlyx7gV2AQdtbG4xRTXkBNJCSc4KxP1J0ylPrkV+KP4ygn10MoWGW/8rR80
bNuwuOVfLlnPdPum091Ejymc+ij2RhORKbIqgtBTPNcCXYLSB7wwb9rg9sZNAPaX
M05ir+cK/bkRtloiTiCNESIEHUVBZHy+b51+4xzlg6Qtt/wxfSaavnTGUvFfYEtd
11YcIfQlEnMSI5+nGoN4QWSvdu4YBAYohosAh/K45BZK930ZC5YljHQTdqLkLXO+
E+VdfgStNwc28vnGSPd98lemavd6DcI0/gRjqy4J0ifdBeovLhaRg80H7fK5ckMl
g+hYO52pfEkf5wunmAi3YKVtn2zDeuPupzHpEETg1CF95bxIsIYtInfKstdE81Y+
5TRV2ka71H6alQ+tXK1g+wiyiMA1rt6gWKK9QGAARm277NgulqKfxpF6lAYdtspN
apaPs6OlH8w0W5GV9htgjD9xBjAB6fBOwwuoF8mBlSANAcemZ4KOigvprJ1tXNCq
5biNsEIKDMGpW07r1UxhEGrpFw5+B1HMd4ksqQydHOH046ALVcC3u9Ll/FmZD8eC
pJC1RC971YJuvgq3SEJkudlW02wxc77xtOBEbWlTNX7Mk+UEzEdP3H6XEymAXOur
IkM0KLxMDk3p8pZ++5HpeJ6JrxdKnHkzqW5YyoqGN4Krxtaq/RRbORocXOn2zeDX
hzkm7CvWVs9baYHiGKzYW8CIzRsPsgIx/+eqnzm4HzK8P9GwItYxWMzWNTOX+Ei1
0a55aJjoVoQFrGx7UvE2gqpain5UpQGGkrp8jNa2IcunG8LkUP6XDB7G0rZuWAgI
Qq2vcXBFw33G1i6zrM38bdSv7jFkinCWNKCjV/j8WLSbwpa1x4vAaTl7O1dK50TH
ykKaTWA4iyxfVK9yEh9MwBafWgwPIqLo+k1hB5Ol76eNpl2ehpAWSALAOr/q74/v
e09zViM9GA55Q6D+9SVBYGSHCGICAHDBd9MmnOK0e01VRCrps1i4HETZsmjJjbp3
ujQJoeoxyNzfhdnqzmtowK46zQ9ipoLDSDdQMspvH84cNRjnuVWfWhQsbUuA+U5k
xZAWI20IIqWlnYFwYq9B+LoTujgyUbpP0efrhtMkYcAG4y3QMjxMc420kyuKBy+f
dgqw8P0282HEf2gSRENVgDYfphvaOiXg+CKlyJIzPEEr/OOGrhy+ouF4IXEUDKwE
wcf7vEgy/ZqlD4wNs6Cpzh4wUwDdFfxzU5eM82A7KRRu4Kp7T38egU6JtHVlCevW
zS15XEcng9zAiAjOY8DVJ0hKoEqfbFUFSnsIMsL5+0W8F+3XyXYvRd3h44C335Nl
N0zpWP4RwE7iEwESRsmBwOK5XJTrQmPjJocPsYc7ySH8DVdHkCHae0TCjQkhJwVj
iGnzAw7VBf62YCd/rSIobKlqWaK6gtsGMQn/xaewmLpOVcfUpudwqhfcIgVOy0/F
kizbHN1NcdVFfhSRTB0EwxcgRiJsQH8G9qoCw8RXIKtIPaXyfgwTEqNdCo8qh+lp
PbGG2kzgamdgWAVhErEd2BgA7A0p7iThNQJJ2pt3sUGkQ96YFGp8P+ydCYdlkPac
jPquMx70+7yMX9jixKEh6TL9bOwYXqFwObqqc/H81Qt/EBv8TRG+NV+xkzEbJ7cE
B1qHtVVAJhlrSxgXREQbXW6rhTCdheWWrQ+xFnDb+4f3Yq3GC1QvBaGmKcggTZGX
XwkACateHNxB7gpqljzomK0c0hsMs663HCpHl9nM1kOWwti64LMxOGSdXxx1+cj2
q2bWvW5bnK6imQLk+IuG0eprqYi5MioC30D1K4WPyNTHc3NWOSvVPUwHheP/fOWM
63HjH5XM5u78sf8BlYR3CqcGoZAuh+p7uqj54BxmdaTB8p+JNQww7y4juToDuoRT
H4xdV+x4xbxkJyjpIqMZaRBnb3yOKAm7MgfY5jDSfMwPoaY4t9dErTEOMRF7xV5q
sTzrzjcfNjxzOm+4OcDWXM7M3BxoAG61ZNdbN8UWkmDT18noRz7zCmMRP1hWASZ4
1sACaMuLuWo5h+QKJhGy5K1HREQKNwgNw8ENc+ME22eDD0879GCOHPRf1dQYnpP9
y9BISSNIY9KfcLLffPO8d4MJbPtg1m7oV2Q+wV9RWqQwmwBqwF0N7AlrCpnVd3eF
vmzrQp+r9zLfp73bvefvQmCeH0DDxFjRItyn79IEpNoE5+m9QZJBcrBxRNW8GtPb
+pa9L8rw17eiG/rqPrDuz4XQRj91IOjN83cyIyahnBSwwa0FYM/9zdsDnkdaDhDa
v640tba6OiP8y8FVq+Yw1i+mBfGFHpRSxwyaaVvOucCV7IexjZzs8wCgnHvIn6El
CGaLTYVhqlT9hMI9j6SNXE3KsfE9tLdI8DPmNKGXvONFZA7+RTbb5g0KbXWQGuA4
`pragma protect end_protected
