// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:55 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
F1+OU7FsT6o2Sq1/ECPquTu49GXbzQNmiRNFxBvBwIqbwk56SnAw8a0Pkrku7lUw
b98b46si3mfp57Fxl578ZlQk5G6K66xsGHmg5yKrYRi2om1m8yG3v01iHhFBQTf1
YTgjj10FMoRfqTXvPCkOJGz2HSgvI9hcB1G7ge1KDWs=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 4288)
kX4bR0POKETNB0R4dLIvowJUM2cORuFs8e0PUkHY6+GDVHNjctrHmaJm2IzEbRou
AKPTdc2U2sc6tGbyFak83mKq1CWGIsIARaD0Gl8s80DjYXRW7YxYJOXUqP56v+oo
EYYztEax/gJgcF1zBoDcph3MN8/gfRLzhLAYO85EbrxddUHzQFYKpJNu3Fax7p/Z
+NAhU3ea9eYeA/FSzWGlQZ/mViXQPSV4O7CLdA7AUx3QjK3OvLjaBATn2l+FOnIn
AE2MuTLKKj03DvMQavpOT6/Xhucmkzu5DpyV/8X2mSt1HVaBiEgebwxxebWJ/8Gh
iiODsWHi8SPicVyOuPiGCnnsOhq8vCVEPAdhcxMF/A/aBwhX2PwUzwQXD+S+xKP8
0/2fkxhD0yBN8p7+Bk0sl9+DHcmkLCAOVmx+s/1IBuXuuhrMsefx+9SXu+4MbVRq
b103Rn13Y8THFxW9mfVx1i3HolOTwJ1S0unw5njk2q1wupxlNfFDVhrl/a5r2VKn
IgzolyufeEgXcPmjq8Dm/oicvUTPtQ+uK0ZBUdIONnYliQDZBD984wo2EIGsqNj2
nCUAdxS9D8zURxHl9NasnJRY1gSsi8yuo0ownjUiIK9cUEzurQ3Eh+b9Hprha/Ty
Qt1X8QeZj5CIAyn0EOANf3p2tDMgxFmhjDPR78vA7+QKVn986AKwnl7D3XM6hFJo
L9UBDI7VtqTcxNHVj6PWzZUupTySDD38MVvgFQ0MmCBMgmZZVo2gwpUaJnllBSGd
Mj2I3C2ziowfbLpTLnhe43LNw9VgAKgz1Qg/0KP9RrzYad6uZ1+MoOK/5A6J9WPq
SAe/EeSKCutwVi3DfyvSW0OVswD/opDpbCat/uhcXRXnW6C9zodw9xFjRPl9htcj
TuVnzmDofkaEI61CTuDXok6vequ4aLEO/HeooESA+DTrQ2LFAWTuwfCRXOVSUFTz
4GkNand5pcFHMtbAAz9ctUjr6oyW5bjXovKF9ruUOy+0zaSQKl8FR5Au6Av7sL1L
FMXkxBFZ1zqW97NdjpY6uQ4rL7EPoImg5tnterH2bsKqcjeFEXh+RVqlO+MIpJMk
nJslryE1NeILNqwir0n93RVkoRL8Hw0zJkx2HtETT9h9EIdZ/ldrRGN5TzND640N
lPq0uKNxrL2fPxp74yIeOaZ+opJ9+pHZ6vK6000MYuqYac13AP/rqezdhhchQfb1
UX2ZgxakbId+DCLTZY9JWyoWKc2daW52ftX9xZ9bM1DQKRFp34OFWu7LNUxEmUNs
Ehi4CwvOZWneTFuTVSLYPoxyaiytvLcTfQarjK4De1R+t6Af5LvL+TQweF5e/9zv
1EoRMk4duF33H4P/X1TwzEB/JSQjR7MErFuQ4iu3Vv4QK/lpEO34QJrurV0dMjym
HRhoCVxjWOlvKaSFesipnIj+13rF0bPl3ZWEZbDvy5uB8PfYXKKqqbE8OOJjS445
gv4GQG5I15s3lwR1b7ONQTFKu6G6TT5J9nab470glVR/nAyYuu/k1U3SihEBt7AH
XALn5T2WsQAhTnE+OTi/LtdOaEdRCajm4SZDWlUlJPUfkU8YKD+Di++aYe90ts2U
mf/pUcUhuKU/lHFQKgj+883NBog6UkFcwQjeR248sp5GJBNb5C1FcHgocmIM1AZI
nYflpI2k1T/3lsmdpwjVWCvUUE5aFGZ6jLwivGt0jJY8WQLYAzTR8gx9ELApQZLq
8CBnTRvvyXIObMOuYg0T/Y3hBkTXcHYu0/FGoy/VN9ohBnTIiI+Jhba8videAFFC
rQ6MMOH31XY/VngsRkClFsZqYsvod3hSEOoEefJQC4jTzzeOOhSPmVpvvvmAOLeF
sq9LIvFGJNxznQys2yTk9etaRF/L8vJ5+EMVsIupBZEhMAi9KnTjml081qsdXnEd
ad2xn8D9z77BIsdGiFshCRhFSbUWHy+6dQu9G+Q7BfxRpNfFdR9prA2Z/LXdX8Ru
Z3fMpMlQRTgVp37F0mDP8Uxe0MT5JfQPUOPl/UYg40Jsf/H6Ovps4EBoFZD80xk5
w2cMoaNlATkDh3PmC/h1WgwciQ60KXgaXaPjZLA6X661BEKVQEqqCwcYLMDB6mNE
/Kc0jylHVLt1FfmwcfEq3ygtjXJoLyHqbY2x1NplzS+NtxpibnhUS03QtxLLyYZa
VlwQ97zruSdLp54W6FRRwIHKWctFVWSv5wOAWGgMIvvb2arBpQFa7CbihrBger88
GnT4voE+3/jIMmaxdz27RVfNzVlQwr/RjyXOk3BvnlfqPEKY0SciXB+sI3l3d9Xp
mcxMGdEM0BsuNhclog7DNe4SJk+RJ0NudaMKb4wWpKkqDzfhWgqKEIJk3FUmXMCU
e/JAlkfy1/oE0jlBS90SV5QFqXKZwcCckiGYWzyFNR2SNwUfhroIyCFv+OkVKsIy
vvpp+matqvJmoAkONFaebIs04xEDyBAxQnTR4svft8x+/FZ7QXeIpWOwQB5qVEQJ
20VWIi9LSkgy17dd4MYIVHTe34ygf47XZvgrN+YnP6OYASYZsyuPqsYa557B2tiQ
0RzcKGAWS7Re8jcSYOn2XoPdakRl8HxIdK451rENeqbXiGLAJGRCxSBATq/1Ua/G
wBGFsZFGtrqA7+9sMyCI78MFQPTcgYFdQLHsJPvsnbpuRgtGEfv0SDyfeuTqEP0j
CwXV3o+8zQwjwk9pXtxk5kiOspd65Gss18nxTUsOaaa4ya0SFVFR2JPxF7aPq/P2
XHZdjYz27uTLY9lrG1C7Tikq6H0QTuJuB6doDDPnE3O0s9qtaB9MbASy9LLhHZmC
4Vu/qqGEAmPXR7Z1LkPrt3h7tNZjqczZZqFYdRNDD87QvU0Ju/XIfyrLMPL2XQHY
WK0Nzmt4Iq7rEzFXbwoJFmCBlgkG5yWSWcaraAARz857J/oPpkGwS+R0GWtAdzwb
stY/XD9LPecw0jSd2Ys1JhsNqlrsR3FdVXb4TxLJLiM58u3lLzfqxKZfgtrUuKFd
Ufzdnf4QLmtqGA7AFCYJ2QwW9Yg3PJBbpsCPbYBHZsx2HmLPVhtSm76RU7QYxw0i
m+kKuGPIDLcnxKwjXDlsTN0q4ZXQO6ZNHwO3jKYN3t65vKQUtBW0OEfus0klm3gu
qPAv6gAEoFvAcrI4XJh1fkTZwHHdBKcJBGcU6KvqYtj/tiAVWoPlVUFsOf1wQBak
AHQ0IOXlO1/qtB3ZgOsypPw1EfDCWeKlSHVZkSij+WrqOMmlETFQD3dkxGOUoHPK
HyN2Ia/PZ800UPiQrAZ7nykpi5VeI2gV1j33lrx3NLmIoHAr9DkRNodp/3uV6zlD
36p73e9RujmIoa0sx1EX6IITbCkPtYJLWgJP/XKMVRx/wH6nnyuXbKxMQtM31TAp
/7lYIGg3IybzYaifX5A2enLgvGnPV4GVw7qxlHpDBf/6IZW4jxW2J9J1grZP0ErR
bn6ME5GelOK82huqhHFeg2p27BM1blbu4Wx7j+zIeK9guWbeVibN7uW8s5XSF2fp
Mj1xXOq+LfUt59/GkAqq0BxUf/P158YkptKHP+izjEMLe8975MBATCia1dygHB9C
3LmeFzf20ZT2KH8fmp6+VVAXOxFjpkIqSAeE7em+Wd8n0pBnpVZYuHOP+PeMW2+Z
B6fHR1oOEn9+oB6npC30PwtS55JhqM4whGV4Mgdorj9bWao6wPA/ZDLi0Rf3w5sS
+wcu3Ha4lvvY5mDbdvp/Yy5fYtTHLqnUz3pt4OKjfxvzGshVwKQBJp1h3Wy1JGEp
pZwR49dGgwtTn4ibaLBF71g8CG+a5Hx4IMYN7CpX0+xlimPPBx9zX2Omo9jVDKSM
btVvGPzU4T/H1Od+8GoNdrOj7zO3vQ7bnysfaSHmGaeDe4VjH7k/ZZ411UFdEXYB
higvWqJoMfYAFAf0MInmnTdxDrtQKFKLE0R6Umd5f2wwJaIGSdYA6JCJs0poSKfa
/9/+Fvdte45cM/EUkl+iZmf7HQ+jKhO5hhV+xJRXmUBPZJeuRm5cCHm/1jhalgV2
a+5Y1VvfAPIRNq+u/6ZAkOsIuFcMwtq1gtO+nWW08aHNEAyDdI59XxgDjUA8VNbr
6pYyfxRL+H/39BwSm8Aarp1zabsIDAnePER+tMK3g1Zzu4/Hlz/TXA3WidAEPXJW
ySa755wNF/0Uwa7I/9bZczNbLtD6vO32OLavcUZJ9mMipGvxKlvb/e+C3+feJx1J
zOS+7A5VfVBL9uAP4pFcmqeHc/zMG1ifwZ4IpNE/LR/agHFCm1Beot7Sp5mJqd8C
50tJ828zTQ14VJ8KZheRcHY7ADeDw2LyZ9bEZwFAF0Tn5ny6aB2qNeS94beDfiXO
nyK41q0ATyIxONBwxRDNj+w1XtVqBr6mGlcOeo5eo3hFVyFJGXD28Kh9Ga0Hs95+
4K0uC0FvZuIN4ziTsxXMw0n2EJo6vkp0uXT8fRvSAAnYtl9mMXWWvYrpz64ZsGkf
nUYCLSZyMwMh0FuXA4EReTuVLGmmaC6QxUJK07Hul/79OVDuAOe9scXbI3/OwzxE
yH2q7gE2kfevX0Lv5XLitvSOgKHVupfafu4FFusrRmHGr/7v0Lbqv/Lkdh0Q/msy
HSqdMPtNQpEtoi6aC7w8nUSEj9phYBgpa/LKA2ZItEYg894n+8mxbi1rU+9rZKOt
jg1z4U/uFWFoL+79WEM6nr155iMcAQ6s66oBtDxE7tC4jL+sIfPOgt3KPQqNQIjS
ooocuCbJpmKlCQH+ZPzi56Kt+Ybp5MBhKwsZcmS/uvH098RVeJGwgxWBGQhyoEob
Ll8sMY2FU3i/ZWEihgpFAYPSNMvVMgG1wC7q+ihCHrjFsNaiVa3YaZ5PToh1OmIf
Qpu9sHGgy1pe+qQNhi7QR6m/NYV7MHwPOA1NVVB0X+4kNuZt+7kyOW4N0HOoADzT
WqcXug4evs/a3zkZHS5APtYiLizKJ8oOTwzI0hbjShBPfl8fvlQEGLTLSlB9Rqva
PtuywJLyIx6zGBjDL0lhirlPZvtDoqKUxmaI+vfRdl/iLVRrEBpbLgJr6c0qOvYu
kV+1rzdUiuzfsrk3vPVCPY8GyP91hSNcJLYNVrtfIAB/b4q+dgkeu8Z4EHkyV5+Q
b3TNLkNGIvPe4Z4SgJKccZC69jJG46vK7dM1+fJqoIl1iSui6l6RPv1rHbl90+yx
KJkyc//P1vcQEILuGIc0BtJ+K6WPl7lGLHuOGtnSGw0w/zH+JfPFOuXO7vPKqa6m
9NhmT8OSLKNT5RjJyqwi50XIRt5ZU/BtHYOOt8Xgd5CBBPu5PvbpcvUUU75Uj+mS
F2dKSRMClLgVcTXWrfFVr5PJJGvnngoV+DRngWoVX5hT4TBXybCIZKqWFsGacscp
83snKg9hOfyHD1yQA11r9cskAlH/Gop2gg5XDNjBxukG3Wq2BGu2kvIfNyeUekee
vZO8hLNXjytWqgMbAx1H5kXWmcywxkOoCghsLxh7Tw+XiypGXMCC+6kpdjn6siZi
v083Tbis/Uin50z3EYE8rzsUXeeTTT/AJqHDjG7h/XJaTY3oIIzoUasWIW+5mws6
Fc9R0j339P50wCjXwmrf67Q2rAhsbyCbzDQK4Q7c4BOtDCylp+cp1j8ZN8kL4N5h
e5KzFUx6FnADlLjuTAd/an8inXCbAgJYYEWZwEYxOI9eYhT7XgFvShpk46BszGyS
kehRsAVmgltLWWbsopBSaw==
`pragma protect end_protected
