// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:38:02 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
EqlMUQmztMguLL8pIGvUGP/UIbzKv+EbUlvKt1eeoWDcPSnniloy2TUrLGDXEGa+
C46HUDZDqloVfhGHOK+E9d8LXAwQHqQyFYneN4X6vNbygpqgUa1mns4BaED56xgZ
4VpBOUV8c5hUZDxFouYxYqHS0YoNhxHtP4tkwyljSEM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 32080)
8cKsTKDvsh0Yzo15cVNrGjcv2iTL6xIAFXQK0E9Tdr9GgRfOxpYrQvn9yEzdzN2p
LvmfVSwWsbhpWTVZwzJYPnUZOImJK11t65Ok62eQOAHX/MlzJuYChZ+rpF2TUMR3
+sFLB218fOoNIJH8dq3oiSjWTvdKOe0gfwpRaPlUEjIiyn/OqX8eVT1POho9z8hn
ZtHCvV/yKtCeI79ZamWtCGy76+QAVNFAd2ZdQMXrFpycjVNPsL7TrsxbaeavKw4i
vRTDgilKSSFjE6V/3W2ZctBvtcKQkaL7pPXTt5wmHiSGjd/PrXWNWylqIBxuLYg+
nJ6pxfmswTXjVSZKT/kvAEjNznr05qf2HIvBE7we+7GlGZXSO6KTYMWajSsWuoPM
C9oyvVhWw7wfEiU3avJHl4g/e93H9IINypCg08p1elNXZ065SHCW7P/K11v/Rn2N
7t2N+TbDl1G4RUbjueTG2v/DDsXsqHi/sEulGwjDvrHeA+KmmWRz2pnnlhhkf6bo
lerANa8DwB+QMQGTBc/lvq1h+wkoHpoKBfYtRz89IpDzpI8TtN+XzcaYgFDanBlT
sSxxKXOvHDI3RMWh9xlP3Up81eRlrdHsGxrohUU4dIdk7nPbkknqwxVpgRDr2VOZ
nD22a99WZADkLfr49cYFywzO0Bmbw+qH4slRiyv4RFiS3WOdwV5grTi5xiEGKlFE
ozWaaILZbo7AOxynP01CQiiAlpdMb01/YN5Qmwk6cFdc29x63ekdGRAxe7aoRLTp
3G2RoVUGaKLKiBuLfTeznShzcFAGsmbBFFZkRkUsfxNk7RiTqoC7uFfVhmY4DiJm
pzyBq+rb9fqx6hcMr5AIcl/afmhVW2gRLmswmQETi8Gdv4R8dAnxYviQKnmEP2Z2
OoUs8eq7zgbxrwoM1bVIdUSor7/nvS68Sm1fIYm6h/WMkpwHx7vT6cn8QXFS66Lc
BlJ77An4O6bLjth+XaTGJqNPm5xkwNcPZgmgPUteEy7C5nc0A7qJKtF6iSaKYItH
FSBz4RAiZG8YOSTTegwL8v27k3tUbEO7sU8hEN5Y+i6QmsnNjpUBUQpVslSme4ZE
UyNgxGH5fzSfnT2WlSfWE5safDme8V4ZurpohOKZq1+8Mv/ZM6ZWMX48VBRLWEIp
LX090NY+COUQT3LvG6PvwATArKm9z/UA5DpEtxmiz4gAp6WfIqCx1/keUO7i5Cz5
g9qhwRky8C2Ck8Fl+NwTghAvpNxVRfiaHIc7Reqc6mi8P7zeIp7gVIW8EUFqaqCj
2BJ5HsCsAAAwMtlM6HflKPok29SX89iLIs+kPORQdLha1gNx6WaXJOetd6zUFOG1
hfnCtgLcUtcBzh2KX4NBlYyCRCm9XIbr/8yZPE3gALPfQtsiLBlLjAxNylWN5hLT
2mrDzpaE0F+vqLlFtDGR44vc/oV2zPFOjTO0gJeQaz7d+tezMbIVmZL0/FkKIduU
6kWMbMJAVr4WINjgiujf66N6zMNnX1OCbhbCMGM/WAC4a7+oN8+VodUZ8Iv1lcZ1
OEgjQRNQBgBp75LPeVrQOqJRHWPdqTuaVGHQCoom17X2xyRoCn/z/5LbUj9WurAT
8QSEsdiRoBn8RUtU857fIjbZ1R0DKrHHk++HewoQZO4bfD5ne9pRtrb9uoV5/wrY
YAHvKp8G7GNjrFqcMt22ZnERNhco+js+UVtd+BoRHSWEv/NOz2Rpq/6ZbzSpzpBc
Js3et9r6lAfkNT1QZaftH10/qWhJhiY4/AXX+BEK/fLPuU4QKRzeM+7uRf8PHipI
HNrJA+vbqOCBWHU9SEvVO6gtqN617B0X89c4fGENI+FHn0aQI/FOefhLvlpas5VK
Y2rTCOc59C8EMtgXzXMDyK/oZescuEmr2YlSPVoYGDaA0xLevdl7EnH1BnxAbUOA
6ngFUpTAVYm/DtMp92rQfjohnA8G7+LzkkO7peLSJYRO4vdla9CL0Jqy+rz9TT7+
P8WRAzCEge+TBxe9iKlQSSsW7vMK0MfTH45jLUFckIXd1JUhNNP4xLffeW6C5Xk7
calzMfpBvCstxv0AZJBGoxPwms1IQxIPdXEgXQ9zb0hFBDFzdBZk1iMQBky1RK1r
7P+OMKGGu460wmkixaxVS3SC8G0X7dUV5rGqfwUdPHh3GXAAi8I8RX4EkaTRVNtR
sSCXf0lnNadguBlcUKygBgDGmx7g0eK2KYfJHUl+x9D5tRXLojPwUCp8uYsaUD/3
DUdydwrwolElIZwYnW0kSQKKCGbI2gOqKT1pVzsKPTFweEkvQkgLWuPOrvVfp1fA
fCnUpCL2JLEkMrZ6h1PBFAFAJUfuksSbSXw4txJXDhv4IVRuHz8c2+SVo13qaItx
OPDpvuw6PjNCH7qdylDhQ/yMfU8T6h9xUEKoWpe5RsBnsahsy19M8YkZfffKfdKH
xcUbzK80gUUHAYg7tfAW8/CZDagG8P7ZWHunjscfq+UqSUgivwUptfqoUVx7PEaJ
j/JemTMzL/yIjgzwd33Bb9TsJKgvuAWV9TzK+z9j8/3e6r+JwI8Jza/HMcmrle9q
VBMRhIPEIm+agenqjnOumcepAGfAwwo0HjOqvve0YuNIa/TI7zQw3ES5sdIwsdqA
pFEZWVp/kdlzyZ3TNukFPjGuwpv/Wa9GjmFMlnhlAKeGtLHd56vex2fTOuh4o+0K
n6iey1SYIhobEkoqp7fIh7KhHe1ewh7FZ6+EWdGv+mI+jaB/SWKnIN993Yc74r9T
fMuYd8okceIggvMTS/6+KnZWUehff9uuizNpJRty6U1KqQ4MSu8I3WpbFrlsYg6E
D1ghTKVyBq+nDvVg+CVFdp3AgX69w0fLVkl048kYTlS6USre4hZvGAPyIrmfH3Oo
wtoMz4GcL9mC7DLVaPxqrHYgJ/cl6J7ehdfJK7ukEOxBqvUR2ZDUn/FsWyx2Ub9w
eo9n2Mjq5GczGm2FasSzptfWiJr2Lu9S3JecuJgyOrjUDLqMWny2ziRMoAJj29zl
Jg4UP+GzaCzzE6N92kBY3gGm8nkI2uxMOfJpNzvLnDN7JNHVxT5BHbXi+IyNLEx0
cejt2D+td0wcnCrdUeyjqah9nN8wZbcgKghwaoGtwQ6Eb8S8slD5iOTSEFxQ+Ngk
trplVeXYkM8HSiOQ8U98OZxD5DOuXopMhnvoXyfcj144DJbgIWF23SZY3kuFC+Wh
izcAzZBGaxwfpD0iWnS9YMKJMc7zmP9Ff4+FLyAi5tjzsOMbQPVMstkdb53ryWOe
AfGw3j1DrE6krnV8n0hFX7zOM3/LTQdxa+WPW/2CefzgagppER/h0ClnqX6Tho1g
pI2o/cRFZB4q0yurX/w+tTmvbYKiD1zssxGpc8E0loFCTLHTMyVocZD4VTaQicy/
lL6lPIY662yPUf/cpBOnHbpNop1VFRLG96w+0G7VElg5w35/243QKBoZLXItDrUQ
N133rCR8eelfvwqILqfNw8MwoGMcHMVb5b0bZ/fAQppDs09E9+HRfGiF02E06dqg
8qFVSYE2T3DXyj7N/fK7Eu8/weMZKdfDeQNMJfKeHbQj+/8kBUUv4j/jWA3Cr0l+
5WjP2znUL0P8dRcgX+EtZoPcSsxmRY6deLAYtnSYb3Y30DfBk9CWwdjSzuqtoSja
adzg/0/ysE5oMVL2ejrjg2ti5vX3ilSOVIvKWRN8Kiv0ZFh5a1JiIMBp96os4UhB
fuouO/AWe9x7NmlydSX/hx+0UhNp/LEciwA0cJ/LPIr0IEPIHJ3qKGLQUBgjB4dM
wSk2r3g9EL5HfBhTcYt5U3nDlvRQbqZX7XnU3HfEeUpSqMIDJvaMG+SWzPaGtER6
zljXq6YHvbXICKl5OptQORJSz0gClk5k7NhYvv7jnDHbVJOzo++LSTv4JWKSEQMW
XfCYztmAw7p1KIzcGNq3H9LwruMnUgkvEowJ+/UpcXl1bqQSCpKedXNOSD10/aTY
wQ/L4Xu59CJEp5AAwXXm63XJwr92yHLXWXoNH9wB+gv28d/WpD1Q8T9Hzcx/9wyG
yzK4w+ItOdxSLblqbSJ4+dao+b4QPgueeXc3NMh45yW/hVCRvcZRRkzt/akj/KsE
R4tzCzTIsNl/P3EUg9a2OQ2skjfIztZ1I0s7IlG3LNr694Znjtfw8H7mBXdTzy2o
7sV+XNiVk31DHpCm5pwrw8K8ovNCJJK1373+bgst2Dml4CQ5vyO05tvOCC/RQ3ra
m680xujeoeE9oYNdmRKSS1Vx8wyQ+X8rRRjflGSPR2k9SLVWkAfqGzksi6YkCc/Y
tkBIx/2Xw4HBWr6mp22LVyRZSlB4YGik4kTb0Q1bzb44MaUJeuCzcYVm7sAhF2gG
gRSQ+3wCXChrd1zL4Y7sF36tQgSSog7tw9T5M4WlO2s2XRfJAWJYop/LkKJraOxB
E7ept/0kSH2pZGY7tP+E4BsrcyEnoOU7PGfA2JheFiNJe4ndOKJeW+OPyv4zxGqr
wCSbbXf1Sa4HvYscbqMLZRP7g/m2vComCdRJ3PgiH9eG7UWlurn/PcOO0raonukM
jyRF8fbGWD8minmTFjZAiOmAWgAAvcBNHsf4e8cFgTOtRkOItMtaD4DehaYDGCDA
1x5k9d/9VRAdF8rGdvShdlZwD90c/8hc4sfL6EIMa013L0imDmflzymsgRid6qrJ
gFkXuhaPnFjqeUoeFN0nblmMUwAUDKVvbVTXDunS9ZEIYH6b4qavsglh0G76mNsr
eSxBvBwHQCwVTIxDK8+itKXjhtpn2M+cl08YAUUwwMR8daue2RuXO9wiczbGJ3Y9
f+LJdBCxwaEQ1B1vsTt+uRKMVceptyv1jnHUw5vH3JKKiguKbejpbiT+J67TdFzn
B/xtjAUbPxoLTtJx0SDGDUZH8vEtB1wHAS7FiD4VyM0XOXKa01boUYJwP1MXc2zy
j//WZfP3Ecj4AgvdYmqCvfIafAwAbDkrPpUkWlmaVIjLzJp22qe+GhQfn7rAYwSN
ucaHHDFssl8OUOUd/RuGpanZKSQJMjj4/WMBpToJ9o41eq1cuUJtjW1gXCoyV5Pm
9v6D+jdZWmvhPwWGOaF5HR6yABC2PYQeYW6fpTx1flN3cU4oLz1CXBxtOEvhtoZB
k9zTM7TdjYniQEN2SIpaTuhVyZ0wM/mQSE5ZlprCEYLijt2cRSoqnUytWIJoUIFx
pHKeQr2tz2gm5ZyY2OFjH8kBaK5wgUhmN5VH4omqk81/zKVPXpn78MCuT9wgCZk9
u/0LBgUjC2Xk/7S1pauN//i6t/iBCutnJn598/ky8rLZi7lDUToB1rONu3biQMCx
QITZ6O0W7Iji5kUF94zW4MmiZTZslYhjSlBmN3qNJseVRIebiC7BIk7Ox4HMEJ/m
p7+BPP9EMkVvhtdQzcJJuDnRzu/ZKChtEm+O6Eumme7zw05paHucYnH+dMm8LoAc
N98qDfnxcA+Ao5knKfq3abaxWEueCbXbEqDHMrvL4GD8k27LVvnKyBt7gXK3YX8V
RUZD7Qw+zx6Jltgookikp85GG2lpHwyOdbbWjKsAv/nR2kLvIKWZs5QMyLnIXcCH
/zw9LZWB/fS19yGC5KrHhMDCW1CRqTMwMpELCbGDCD3zsKcSsXdrve/CLHNVIowE
qtutt/hdCGT+0qzo2yJMvEm6GXLpnXF4rBK0QVyfLmPf+84sKZ7qVRlm8sTWbeBY
HLRS8puy9TesLu63+RJ0EqdGsrt3O/6Pwp8Hf2fRLMsrnzRj3pP+X0iJIJHri/XL
N/ifYioNcA+bA4ppBOJAgNAyTL9dWErac6vsnBS/KfS9kmMPiJUcglH68DY8amDB
0E35ljybEvmVn9m5Yf3rjM0o/jCS9d0Y3f+6ENP9G+hi6Nwtayhc6n5VtxNUeL/S
daksbSDLiqD9hQ+wjkeHFbqJIaZI5PWplsSj3sK0l55J/dIK5XyzDX1x24G5SHvL
TZzTXgIQVzQBT17NkCZQazYs1JQdlzDN+RLqSJB5RSqmUEbj7t2qhw/X6uA41bAH
zHswWHOrx1KmcXbxX0dGcb/IADBuS+8Hx/7NUYK2g2U3gxJkiPyJswr+doEm9Umv
+0DUDn3AdQQQyDoF/LDgo8f1oBQ24tRQwPURBbKgN2VdcT/zNQuYeRBkDIM14J6Q
sk6bAG+YVYE3ceYpvHPTxbjZK+xGrk9mhpdq5+beAb4Iq2T95T4vS8PIbo527fDM
KHY3WlbTl7qcHgmpqHR41lrY4X1H/t5t8yzOX36A1nLdFxvbfWgkp/rjOhA9YyUo
iWD186lTMK5fkbVLcdtXS9ExgmOch2r34mhC20F/bnZaxDePE2Iqsa5AQCSV+kgw
NO6mdBDPDFAX+ztpZNsgzCBVqQoBtB8jJiH0GRx69YJeCTyD3D7YG2028ca4ZQuk
LwwrdWZJIUYH6CUuQsEJZhWlC9yWRRd6QBM8/gswU0BkhhKBgcGvWgue312VbDwP
02nhZZVqSSY4Ekbm47c4XrdDZmkOhnuKpgpYKhyRq2lCb5xlqzpid0ficYLfZ02r
0/2r0UbHuznYB2L2G/vRaj1R1bg97Hd+MIc87eLufFUa7p74zhfChjmctCp6itTW
keONJCBOGBukoxCO7glgkLFbJcFliKUvVaeXh/+3+/QnWF5FBWR9vzqV3ujDTTar
t3rGd8hifTX0TOn1/AQjZ6DwszG4mUpW53xQU37g7j8QXejIh8HadnwS1oQiv6rj
CpOj8+HV+FUOdMb1FvstHC9M1GVtqIITehjO08G2z05dCGbQJnEsshqDBN4FjNKH
V/7fTC/r36mlU/xtgdd1yexmCQ/ECcLbv6kkqu7E4UrFGATwQe2a5vDtZa93AV/I
taYt41s30x9wzjHnBXYR+R/eNhvOuBtfNsfp6gM8ahsBFg3Nfgec7Jvp3a2Imh1Z
PBUdmvqGEHV/WRIzVVyGgdayfYZ2a74WHD5oSP5BF1cDnYMnqIyhepHenHlrH4J1
kyHMM4R0nCsIJKb38A8GAfHSdrYeDRrizB3NcptvvFbk/5zX5AAltgTcI993QV8Q
ZpDj6VQtJQVKmqudtJxJLdDLSUXioCmiHb3XhYC/6UvCDXOU89ihFHY24W7M/lZC
MHxg8Uow+rYswEYVRrlJidbDbecqY8qXv/xuvxf3lqySHZ5UM7P7Vg+B/ItHuClk
PPDuzmXDWREzmPDJ7gwUtDBK75FnxNPAJv0Nsv+bsQAzQnps5sK8E6p+6pbVEDHK
dMCMjPMPTv/VjlFnRN0Io7sYC8YCpBRNXKHhl9GxS7RLcXHKoF2tKY2xq0cl4JoN
ACtgQPOxztF7A4DeZOShfgGNR8bZxFaVyaexIH/nqNxztAAMRY1z0ibE4rRdX+eI
0gUiDmS9o0eJAwuEKCQN7U/JxvSSco3wjYAP5W7QBqsaOLnqEQFJp620TumXN2qL
pBejLAn9EZ7uKWE+gVT+e349CPovoJDdeez78dYyfFbPMqQrh8truCqbQaq/16Tc
HhPV1eLwgdd5yKeBgWnJdrdkk1pcV4GchLPXIam62vJIwTYFyAZDrdPzBD6DddwU
9QQxBCpNtGHPoVYztS8BHWX+uHNFUBI4lH4XszRbh67h1Iq/i5x2amVP4z0eWcv8
0b4WB2OSUkng3TuExg09eHwvHbJvGY1PefUbocI1HjX+LANpxZ/fJbeZnIrJyBET
4DKhtGC4rY90nyYZy+aVq3w1ekXfVoMpj9OMdIb3b4akU2zM/bWYiAZPFbALKaO0
gpUsZ63Cv0B4YaPHLG/8CvnzcptC/q893elNHq3TnjhX8y/mvVFGHuRJJKsyI88T
bqv1GQToywx64THcaDA9GMv4uj31jKBruaZqwmaEbnZE3yXTyd3ElxmW9txyo5ha
pguy+6k3G8rg6Q4LIIhf1HnKm3uvzbbSVg8l39Ho0gUM5uDOQxV6cs1AthXletrZ
QbowtAqYbSshKyaAJl9snfru+qlz3VKTF88H3MGmpx6X2epSlSw/6qnVpWCC8k99
mE7acUwoQGTsX4Iidp5Z/O2HrguhiN1OSHRuh/24jKG0hv1rTBgy5jxYFXcuydjh
6gHIXCQOiwAWXp3U8gTlrVKgbkNSgX8tORUUGnaWmo4BTcl2dnYTm/oWrUNON4Jg
D45MV6HwMf/V0ISCXag//z1QB6kxr1hYRsEjYLpy5I7YMl9P5m9hMIZy8bKJpuUl
k4IUnBAFXLxePdnBEwzNWuhWF/CDSvmIbFZXf5g9F6MyYQfgekdRDiZwkuPzvZsd
d9m09RQzIYczCxXH5HmRTBpr6c5KSPp626L9C/E7vzqEU3v2anBf5BW1u0PhXSjJ
Ru9MpV/JWRmM+fjljwL1QYtLkZIiXeUSn586EXZtzl8PdbHVEFubA44veP8xMLff
OrMNlHRLInN3kQVBWmPNpOX9XF/qBLm8iZiPl0Fr8ZuAYgYD6Vqq+k8JAAZ3zCFS
+l/JBJGnQhx1w7D2VqLfFWphmenK1/Mwr4RaQOtXEnMUzzNlYZitQh7rLRcg2UdA
mswI4/bI3s5UE7eBQqGNNtZXNfdwC0QeY6n4XiL8E3daEEPHb383y6QvSQo0/opE
QV+P3OJTlXMnxWfx6o8nV8iAxxPo8XlLft1q9IthX6vMo7rZg1UELdLaAk72rVt+
MzCZacWK8qHMZ0NdmaqETasI/iOpjuoz04D0ZXnwjuWEPK6ocOCCypnESEZutc/K
wb8bZ5f/p+hMWV8b515d4zqJ2ImUdJPDE+/68k17Qy2nwnTMvZiRgkThITi1CD/j
KFyMT8CaCSzuxTP9lgwihZjr2SW+sTxyHDhjiXK84bk8cIQFRUl75+g3mVES1KOy
E3bnAswRCvYMIy5Qo94NKLkNX1BbXlzV8ZIdPkErlrL77clC7JJg6IANghxGbXkN
fBvHDgcc4/Ry/seKyxo894XHEmX3uedaNwGGyJMdFsI49+Goa7G0AY/+mR4gH0lc
W/wfFL3PV/25MJPrcBKhk3VnRqIWxoGZJXiuAjo9avEnBgDl1SRQ/mC/Zn1pRqk7
Kpa1Xd0PItNnu5btsc83fsNj11gp3CI0ys6zMoTjh1VLfImyWe0JXQbBz0+zxLbv
UBnUNJYWkoePVp3JQPeLnOu3I1tbrWZplYQDTpaJ5qCmkSrcDkmiVr4Ds9YtR6xo
bsvIqBn7OW/F4uFxk6y/bM7G5sd2v03ieL3J6cU6o1nMVIWdY4vskLjAy6/h00dd
fu0oTJy9qS4KCPB+jA7dooFq7YpJBKgm4gM5VqpZOYQPYim2BIgvLmfj8RZFNPHr
5MqxC8ybavZ1gpu8Lg/PpV5B27x4W8JD+wy8rdu6v9NcyZINGbDhpvLoUlEjTkvP
7ha636QaaUBgfZy67ocmBMidFVohXGP52RWDLrmsbMK0ZDTAJDYrgvemCuE2pZ2V
eea/KQVMM851JjFimhQA8rBWan3VoXQ5G6qBvmPLVy2CrMArEpkr4G8dLWg8lSPc
ZZzEhgJ7lHKrIsfVWHYTOha13mEoDAL2xakigqxbKNF+aqUNzyFzEc9zUPzbfrBl
Mt0o4uZIKe8/4FjG/nN10jECSvi/6p1YhhiZNZCkdkMfumCiQhrjE74h5FGbIvGm
/lL6E/bTOu3kpBilLthNdv9B7BIbbaKjHicCaqh/iljd8+sjNxsz5TuX6Z6YVzlr
gz8xTlsYcw+fgLMOlmkqlj90fqf7v3He87EmU+rgfBqJgl0bmLDY8O7qcw2EZfWF
c7LhQR8AB1a8Yhuyjq79J2bE0jBkwtsxKANCwZPKwmK32AO8Aq7xXEEM7eXwhPJl
E8JI1xzUCweY3VXWBJ16UcKAgGjzzwfAOk8igEOVlXlvpUqrUh6ukaioi8NyOX5S
ywhhfaoknsW3VAGw7LDv3u5pPg/d+PQVqCjFoLJWDSyGJSCZoqylgkmNseFSpwnb
jSEL4lJSyXPgCqlt8zTwXNUb5WVt+iszucYY+niU5g+46J4Hv5THVR3+nGy8vTMD
ljMCZc54pzaUZhddjgVHxsLv8ndrjRR49tt3GELdb2+oTtw/rgPXXaL8eaAPY+rV
vV/KiG+QSFmZ9S4YKthO95fc7KwanIWea2EwOIzoRw7XaC6vVPRVCwwacQROxjMb
+jMwFN5XTO4gHluFZFFkpoPFpgD7eWmV0kxxCdzZnBybiqsH0WWsIn5lq333sEpu
nYfS2m8/pt3t9flbgkQ91wHFu+t7liZSnAbJn+PzEDadAol4K6oxOkNxKJFYAD2k
p1KHuX4E2Ykyst7m65VTRVeDamngoFOSKrZ35MAhtJL5o7ym/RWdRNz+noP5N0g0
1glRkRuPqnylgmnKXY9ekp7CBXzdorqfE2O39GjFXLJiUlequQxFtqb4+iBkVXcC
SiiKQO9c66U96lS6jWMAvJXMSoEvt8f/kpZSJX1qcEGfUFStKYyZVY13FVIB4bVm
mhPFS2H+MgMvAcHGyDf3gB1BS8EPBAcPFoLT4TGNYlxhhqQluMBhQUQRNJ5MEI1+
iZrZVgUf8sf3SmGrEq7ph9P6hqAlJ7+tV9HPzC3ZiHyLNz3HPc1C5l646q/Iaxsp
ID7JkFCS2PjYFDdoBJc4CvJGD8wUrYXoiZFtWQaPrtOL7JYXxT7l8wCzKSqwq9P/
wB/fEfwjR4wFjb3AhFsy0xig9qdE3XZtZp741PGZHHlhatAX2aNp0kFQ4BYpqyX+
mHuxtdHWnzgRu+Rp9dk+b7VHePptiC2raghihyWqAce9P+r8V+0MM3mlMXL5VAHS
KPZOVrvJlMMMt7+zg/HxGUI/I4I0AsFVLzXlI0TuF4wHT/Sdt8tRTDEEzgjYrNCO
elE0hU733l22wB0Nr8rSNxf4c8MRDwMSx5hbN3Jb13YUjyK10sUFZfA2z5KnovJ2
xDakllXDjbFU9kAnAfM/sETkAK7jwxGm5KrGFdf6TFm35m3WLmVNbV0Co/NKoZm2
dXaFzw8SEiUpUginx6lTiupr2+Kbr89qdTjAMx9HMfoYY7OCms34ZwVzqxlCAVJx
GAvqCUvDVRrA8uPiHErjvDxzhCLhRhx0qBevVDKPezqXuq9FmS/ZMO6pjlLjRMkC
edNOnO1l2WrwXtM5pHaEIeaKyvzwU1E7soUU3roLxnaMugL95rFVWGjXSxVO/S2m
LvdIJN1iaTYjlG9MTT8zoUbO7eNroUDHZ2rR6hZBTwOqQ5ivhDo9tedq2nd0YD4v
7uE5niTNqHKq3uavpiwY5MaeyZoas5oyqpCPHQcWvrGhmMm0171J9EmBfj2psp78
v0IFiGv1UnyA8yjCY/eKWOMBH8VZcLzQRC2T9CnGBsSFisNPuYLUwps5CX7k4jrI
K/A/S5HU0WRDiikvTrgcZRSPRWz9y/Qc/11bWWl5YeC16OLfL6BhqkwcptWCC9Yd
ynxxxoccHq9q/XzUcziLNRHKL4HQGHFhPL12GPtYHjy1XWzTzGwXt3z09Izvu1YI
mrgbnNumwF/1uyVGkHsEC647OaWY/uPEIH0wc+slZA4DssiZ3+ALAmv2Xw+MDypO
OfOv+Sg561CZeu5tuJY1ukmnHDtZq8t1fKbvCtvQPO9N9Z/X/L6yeSo/dPL0iITz
KStZE62k+J3bPzQvIZK1tlzI+jzUB5iDA49a20sxm/UD3u7+FXmxoeGUvSVcFSPY
FeN9Ju9IYQfTVkshBBYg5AhALgaENRC+4TtO6ogT58LROT6ftnCMImdFJWacUH6W
sfMbmewB8BqK2T0+P1/gZ53JDDG99OUx6xGzNnHa/eQbm9kJHGAjzKEIt/JoDWZy
7SOrW5aFvnJOUrQChOnEb+MCxxv2xECUwHqjo/uPApBd7OePYfFftUjcbYcHnPvM
if90cRIFq+mSY4swsaX3MaiaWOhJWqzrY3XF1Y3+cGIWvU78TJnfneVvhxuLrSij
PAL4zJ5AdkWiXcivSv/HWGD3+YlLnyCFWHlXzeSH6a6bItbuXpJM04Ffbz+rZ9j8
cnvMK2YUQ0DiNMVAr4m/F6MnF7bZPsyqhW60LH8VSgdhT7jOeU0Pvkui+aB0vRyo
YVyxvh24vRwrIBnB0R0p1Ll3pXxKXTnRl3CtmLTP7Q0VzwnEbOC1gIBrnqKUHiWM
mN5bRgxV6h9dXMJgRtksOQ4nEYTmAFOXZVIiFvjgP11YZCTb0Qi7xTRiCjnmN5a/
hIA+GUNIgoQE1d0kETyzf+hvSsXf4jT3i50l742CvtaQSsP7nVwnZKXR+ATmaOWQ
a8P1V5APav9QBX7md3Z8a96HWiX5Sc/dP9IrCW52xXcQ5hfNLsml02LpExB0BHDI
x5lBA+Rf62mg5+sj1/y8TeIQnFEf7skUhwCn5WLiTm30beC717t8HV233ExNWmTc
wOqD1fGmgQKt0OhcjSpBzEQ/PgutKoUZJ2FUQ1of/tTAXg+zC3jH+OtCPKxxsUj2
PdHXRy7DF4TYLrwDDZfvns+/FOVb7krKhpxe0tly3DnTUWuJ/tyGBkDnPu76qsBj
bJhPX2HA6B7lBeFTBjl+Rx7n+gRd0HqFFNgVevnwXdu8pXtjfF29FzeAwvS8TAhg
b+XSztn3eOK47GU9in7beyInfnpdO5xpedUWC2iSNhqeAcxpFFdukvnALBFT5x+E
1GJM24YCNkCuoe3RWRwVsqw7+iaphAEQ7vuuBWoczYdXe5S9uvOntbALQXznIdct
r8gGqVfSs76C711jipEQOhnkBlbHI5ttd7es1f2unZCYbXquuXIUkHFLcVMvv5e8
7+9/cIw/FR6KiXcuOv5fNK01DkFB2GbxsAFn4Ubkwrik+NX140W3P9QzHmf97CFT
dIqS69AmSGb1bBu4IUWIYnkc65ctVOTNq6qMxkYRg0yRKTUIfuSEA/WZuy3RT696
GS+lZd755sPbQDE9iXG5RVPRXr/fC4kR53uqAoXozx8PNtJzaj7J2aVLyJ8n2YXE
ktBXmL6Yq1LREygEzIXjIIa0nFJrcYlDZVBpb6LyLF3sZ+4o7htCk2clrviXCBnb
9SCrjXCOvyVJ+9D60pXCNf6aUor2MeXdrQPgrptzgHl0AGwkLTTwfsk+rd9jQTvx
F6BH9GiHezAbxC5VAoB0NsUaF4FseHI856s/p0BzHpf1XUaepqXakkMOKLf1irpd
HEuVimpfAHwZQq9VdjAH+KpKGZ2m2Nu0uyXsOXiN0PA9thQjyQ4IcQY2XlZ8fZAR
8FmrNvGqDoL1cBW4jFHtLa4BHio+Dri5SUFsKZrtLWeBauCcgCgDnY74QxTPZXHH
K3vFiHcaxu9uoAX6gdBvOfBT/8LcVKSu0m40w2JAWjrDnXWDNasH68ZXAGzUCDOb
7uayvQzDsz8sRkiejIj35bVxtl/6yaauUUU8IpKxmweBxxr29NGBvgfqABLUtlgX
Gt+un7yqbpQOaHqK7fw4xej/eWFh6vfdyocDoFyxUWM9+VdbwquwGp4inoV+SW5L
fapBf2h/CzIYtch+UZ6kQ2Ua9ajt7MR/HBAo55OKfiTejz7HSjf6G/jzw5VH004S
UB8j+083Mgl8Bjjsze1jkANW0ubZ5YMf7kaqvrdh7qrMycEsuz+vMlvb10OhGd9B
R4T3FEc3MkwiEYrSfcvpyPLt97hfrL8uHJArPEAfV89NDxqhDbgH1Rkmq8Vg3G+Y
1uN0n4MKwJ3Ap/4hH1XfppwcJogWGtHKLUwWuVFfJ+3EIxOrv0PY4mkXXToYKFqR
ZwnSmGZU/2ezWpMS9hPysf7Gly7olhqfzAWfEcn5soPWQfa16ahR8vyyfRzAVDQE
ds3zfSiY0sru0yExyNMWlXrfxCezpF3PC29fbKJc+WMTSlMAUy9K0vPt6rQbffrc
aJydyPsSdy1hjvH2jIDmDP4LN5nY5a8PSlNngJ1hE3Xxxuvr0JP5Fr0ngHYUF/mN
vIyeOm7rC+dLPbv3beODWZQ5kxp3Dau+hFxgRW5zVX3JJL4Uh3S9hAYQqgk68xEW
VFb2pSEcNM52g3DKB8HlsopI4PFEv0IIQdOelRgvIqvITlM49wX892cOcz/v7wMK
dwRMJt5X7OJcefJGfE4i9qOOBVxOaWVNuAzDlcSa0gcIJhG6m90eHx9J/H1T5aHz
aV4DYy31LtNN/2GdIG5a0DdXaTRjZ03vL4lfU5iKzcZ1bubgNQb11L6GiGVBEQGX
3cfUOcRbmKbFrHbJzezUj3jcxuMJePDr44K0Luj5KQbnQs5VhkWY3qCodB+2ZA7a
kqNOgFThj6kNAy0KiqN4h/jSHwDv2It7EMZen1P58gphFMFFOC8wsFuOJXIAWRj+
wyv4nSwHlZQaTY1FX/JIAIVN0p31bDVUdzcOcM/MTIyzoMPp9KD4RFSnzvXASrVj
syz0twbyNxLmLPGcm/KP8wIMJwbzauMcIkj/bYSH4N1bJ9aopjuWahErlyTxMB25
lv+tB2l/uTyRskvKeMhzaPSNZDb4WkQ7M0vI3upFs+9owtw1XbV5daBfUl8A4SZs
/Ak3n2AMPiofG5HSy9CchT/La/8UApUOikvAjp92ZAMheUQybh5Fte1NyCD9LcJY
OUHX7ez2/cDNcHTZIgrmlNIIH+TyCy3SBLWSp5vZBJVlhUUK5caCPRgU+9pBsAuz
6ggDWv9pEzY/POCLhicev8bzcWwjbpV8ESMtHMRs6MP72I0GSg6EDZvJ1U+nYWcd
cjEDfiTHhA5/6+0ukuDXlVcgUR4Yhaba2JeWmgtiwB9iJx8vwBYMS+Ru3KcO0m0b
Lg2xv4yz08t62C5N8DMtGbXipHPLhxj0B/cYD+RTwU5LCHwFYPEVI1FAiOnTq1pp
BAY5OBnrIgm+VSWYJeOUf9dyy1nq+nQv8zwWqEwonH3uFGeNwni8eyB5wSlyq5Ax
WDXSCSuM+k9Ozc2Mrj1lTTQ5ud61OLp+fzG5OT5aT/5Bw8/NPJc5ZYCcusD9+bQE
BRKtsLiV51kxB8u218mdIZtvHdBOEN+1wBzNvr1E1rLPNnrSaM1e41tWwuazCsBQ
X2iCQ5fu8RTGDwHNXZswOz7tCIbuspM15Rd5RfM56Qy8g4HhwQfOUEG6dceJGqbF
WsCFjIPI9/WKhogCOa3Jwijq63ky9uYmDsPgqx4irnRmevi1Nx0PCAHHgVi3qLGQ
eTHBb9/797dtpXuvzbbhex6Zz1Q/BVJEK6PaDfGvg8+SjwMF1zRoZ6TuFQvt2iTI
ACH1y+oeknSsty0Vk5CbiqhDhZyQXFxq1EolKd6FDtAn95URnWCwW7mp1sBk7pks
ItrZZR+NTKQx+kxKthsx5XTCct8bHMpMVs5wEFJEjsv37UBpaThfBDbi42bUJa+h
jtkS6rPB+/oMY9gD2YvbLolG5qg4IJ7OmujKpx4Guy7vrHISp5La13RbzbxskQFk
BhHAipolZOMzbmXJuaTA7zKZ12qXWCS5B51AaZpxqYWX59KzCkfpezcAJc6WZhwY
RarIdF8RzIsgyCE2E8pbCreBhOExiVX/33eMax+rNFYJPxt/Uw90c3q8w8dfcgev
yI5eoZJOj1UE1R8eQylQlurGbpXtzNJianYJs13Aj1TOFyH8Oo/MENOw3wXDsQoy
PcPefMB4F6cO7QsCcKZ/+tsEuP/8eeLvGTwKWFBLfY6RRWPt+BzrDQXaXXDe1C6E
2cWcQHX03sDqkUkPSt6R0pc6ndsywM0ZPDsvK9a1DRTV4fL7o5ZRkRAzWm5IjnF3
ZPEOhLbhZglUL/HXDCURC669xL6OMaocyOnMNCNl8H/nnks1hwHeTYt1uoP7AFUE
opVdsg8EM5VB0FY/HrvGuNTjkZrkwTA71gq1U3W2+ooJHT4bQjagEM27LqO/XfaT
2zw7FRgefMAGTjV+qbqNS3T+Sn2lAnwiOtUpcRGZu7kaGq21cogBbNAn/Is2hoRp
C/4OhJHo1pALCVej9LWMLqqzNSFsQ2D1+wTLQ+r2iEVOZJGZazMV+BPU6ggFhmSl
xHNHdfNHJFwiNRTGjF0G8k4QYjYIVvsNENLUhr51BQZl35Cv6EO04nnIzSjBBEPj
JPbmFFyJC6tin8Jz7K73+GL1Pxj5uU7e3n/xcr2xpK9O6joJBsSTWcWwSnZTaXpl
VIMYmPHJO8qDh3JzwiXQSdrERtkbo01Bhwt3v/OlUpR1Y79Slc2jXB/owq6gxALa
jY9KuKJF/TPNEOIAvH2u3/rf8x8PXt35tnAc4lH2+sLbYVwmqHq9INboxa2HsKkh
TsVqY/3IVhF5gkjYY7hk49DceJn7lyERYBmNpR42DAcuZUXv/31pgj2CWvO3abcB
y8/BIa9jXqIQWTdWnljN0PEy4TIsVzge7QSyKPKjKIFka0Cg/9RTTDC6VhF+BIUl
9TQ1+Xl3O800xaEJOtdtmhy3rjXJ0G+P5iAmccmonDKgDXsTfipZ0lULTL9Abq3K
X8M2SdrLyUFyMowje1qc0mfCJd0xnnEq9FKx+VNXW1tDqPd/ae8fErLQJeMKWeBX
SlUkrid8tdc/w7ygM7DhcmAyJHxgYyHRpb2/Q0STTeD3ne24tm96lpquPd04jU08
CG10KIhHXGH/oWbukf+jKat+O+2dEnGMhQ8k97jxfHyl9ZjHCYyhLtsbPH0vKwSe
6v0JWouUkPawmx96jPdGAYvmQROglx/QsWHfFutBKkrJg402B/FgCY2G95qo4RBp
0RrYrOy5DlJfDFdsfb80iVqxHOsUA/WTyJ3XblTjcJFArSnbzqZxrgtKwjnJm+yq
cJnLY168XD16iX3R14fc5fPzBCr2qRb9zDqlWekGES8+QDrnvsLB0FQgs7te+aVS
Gitx+Rt2rq66kODSBDWBTbRoQnXIK/y2LcXGy8fQ+m/jtceNV31uc7p4VQt+nSKG
3nuOEBP1kbA2EEMsJbZUmPsA2z4cl8JOBLwYuSULKC6eIv8yPUB2+JXpCLV7ah9U
+5nx274kzPZdct/05JeMKHmi8CxK1qIrAZH8frOxaOFt9UpKRr8uJv3LujRiCrtz
A5zLY8tIthRNXXzyyUZZylavM0IMEqQB38LTDBB1Dw5WRgwQC95YVdPqxRLgiti4
k3rhdHajyFyZhOb3slKm0IgFdIO/lq9iukZSqSqnqp9TdYeoXmPxRiNvC388p+Ar
6zg/sV5wVDXJG7/HSy09ERiDqr/w2Og/VtYjcZ/5yPT1lFXUBenowfuey9vAnkn0
SFi6Nc0Q7Swc8NYtR34NqGI4rOAnLiB5lRufsHZqyTs85le7ZmQlHSHxd3HQrgOu
hjYss0AhAvdGrEbJcIp+8Lsxb1HQwtHbW3bqJ68akYqQ57jMwkybOTPRShagcSqw
MoN6Jdq/t1MxTavD2GW92Cv6iTJuE8geunEVmvV7oJwsarSrmIAoDjNT4aycl3lV
Txh8/Cy44kv3T9ixy63ZbS03A4UIdQnZSgDUrACnlsWQYKF8csn5JbPPHuSWWbQk
INvMFytqzo6nyuha0BKMJ42qFX1/bXmiVGzbXHfuPX4kWAm3ES0Di5b6WKynrL0I
vqruS2cPNNyrU5AKaNnmG2BpnHsiIbV+A8RXyGTueB+rCmicGhofhAPaL72+HbcH
cY5QNEH88nQknJ9WJE8w9ROzlpsDDzPLDdU1AEysNbcKKNjtwAuAkxTD1CIyUOSd
F6V3sZ4p7wDsQq7yDdXTPXZec1X24y8NqeF5yhvp9F98ZaSUd/8Ciw+l9HjusgX1
RBKOm6JgKGnqEkh8PZSlT9JMtBzg2I8jaQv4U/n4ebPDRQnpDWBbBQRtHsi3IFCa
fzsOueHviXF2zJEV1hphTApiU3YC6jp4EqNW27UC0wQzceNcGNDNPa63HqbmI9OW
mkupY2sMPtG58P4ZWrEg5PKhw4i4yLj51Jd/ByBVU7FqbxFqBHmNYvwXvfdLKyPP
S4p5V60+onXj1fgjtgDuG5fuSrEq88MBb/Aub1Z9DnmA13RNhWDbsIjcKEry5ji1
OAZxm6kGVrgeHj+F9cXap3GLqEfisa3uVQoxBCPZ5zrWinUOmRFqVUZlcU4KhtWP
oit6/RYkAzZsJPXFJRK7rpwJtEN70Ll9bFTOMzkacq19725xLax3BXnUn/Joel+K
+mEKvc+3nanB7HdJMI25zItgDuh/4toFWaHZnvPvDrPHiLpqKZIH9QPFSOhEg+oz
r2IXs4F3Gl7pnNFTyfsH0Ht00HuqvN9IAUQfUDZ3O2BhaaogaJWh2hJsaoxvcuiX
FIF0h0FNU5aBLOdUtK8RSuvdRwmfpndxDLMyyzZHsyFGe5ErbSxx7alelHoKXMnq
XHYZR6E7LUH6WdIQVs9Y/DNFh8i89KkMdu3HAgmjMWQZC6DofB6/T6xCvegHp0tV
YGRqBDSUI4+mOxOpKUE8iwl+LggGYnykTg4TDtQ2wjCLjg9LbMbiWN5sqMRd4+Yr
im0Cs2Qb61sA8TwpDZ6IiTePVA/fj2FyUFIfrMiMezoQwlWXhACqCgwRJygpA2tN
CjHaSLF58quZPG33vIcffaK5IO+YjbQ7MwkjUZwBwmL9TL+2wG/actWAyal1YzxX
HykFF2Tt6BpTvLIvzJOS6gjvyLlGr5laFCoK7xjcnE7AK0ffHJikzAvkaoBYz0RU
q3aplrel/6QMzWFNYi5DfGIKpa0tHPgS8lGVrjTLJx5/fSPIugbsPHV/UfIXsvl5
wrWxQ2Z1OoQircNSXMCF8ThAN1Wln93WHCFnYXvGuF6LNYeFZVcFFPujUIZKjJJl
6f/90MIxyV7BoyddfIq0q+UT9pAp1YXTIJVg8SebPxDm0lmlSAYYNwjMxVN4F129
AKzyw69YFRegA4p0Ti9P/hPM7LNW4b/nDjtGviA2Lq4hlSdpyFDEv3+wHtebmo2N
hBGN2CaWPnuqe1hVWuC8BaSpLmHIMduJt6byekEBoVVw09Q6aZXGxs7BXJfROfeO
CrFNnFom4UOvPB3KH+YqH2UYQAImDwsNmYjhEDVMNL5ofHUXA/OwdZAaUDIS86pk
va7QRH5eLrIVTdlnl8rhVioO5jjDp+7TfGoGtnaVrwqahi5vsdAZOq1J3GEn1x/v
GJSfmxv+FSwsqXW8eKyhS8VAQU91xTU4I5EVEIwVsGKrwf/jdLpbqjwNEu9d6z1W
a5K7+bDbkn28VdwOIaQq2NdNT6xKLqFWJhTA22ZuZ1RJD7s427jfNS0pt1qj/AN/
oFTs+FC0LUNpHHP+QCP8EyzneAAlqod+7oiy7UPBUBa4TUImr0lOC//yV1cx1wqA
Gv7Y5qKBqO3/Cy1Nm7UO++RYWaIVzl1yyBTm+pQylkHP6nmwa/dqXySw2cojO9Lh
k2xQdQq0i1pAXfA5HPs3T76/M1uTPk/BqjawawckbwLKypJKBCIy4w1GKoLLy5ZO
6whzfMG3Dz0u9fWSy+av13jFoL01jCuXkccDaGnPBhhvlLIg84dvN5ow5srhnzbB
SS+4wz0Rn++3CMn+LaHv4GziVarq16PTnRpWCelYmX+EiZY+MWgQcyzKFjbQy/hW
yV262L58dDo+j63exYoqSJNyATZIaeQTFhFPbzgJcZFGZvzpsXAQJ0/PFOW9JVjt
9TLDiI5rFfNsDVt3V9B3W1+USGJ1rPvhcjTPvzsfrciwmojiagi8xK8tRrkofOQV
fPRi7qQUUMHzhAI75deMbLOEuhuW/ovrS0Up6dcIHK1MBA/RMpCOS7UnvzxH1yup
0qQlZv+Mk4dfYUNOOC43L8yKKrr4UrrkmEbcz4fEBlC2b8HMlkJ5lvZ0phzqLuHD
S9AgL1ud3aUsUq9147ye1esSwxwma4A9zR3ogBSfUtErsxR3LNGD3QnzVh2Ow+SB
e0iiYHMSY9mWW7txbJstcZXHCcySdfbh/nSOSRutvwrdyxYVwXdcEIl3NdAyLXhx
c6ZM1/5eDTmMI1qG/+dAUZlxPlpvBFzByCsajfUiuPqEQAQFLUB+EUB4F0aKQj/L
2RgTHYtTYMHZwnOar7B8QmO8aFUkVS3h9KHzriGooH0W0xDrcw4F4Y9wOVsTk4Of
LFfHp0/XMzG6TYeY6wAVfybKKHp6ZfDYJxGY3nUc5HkTDDA6ROsa1bfChd+QCflY
5LixFTeaoXmo5ho3EPdvtFI0JUetz2eEi09pgSUbRsi0HQ1/pqRMx555klhHeOHg
Em/6sON+UzUR/0S7WFt0zExBSH6sONlVyyNuj/IWehRhpU8bHgM029u9PNTyOr/K
54XWEXfj2wAk49A2q8qY2EMml1zX0yBnqdPlEG9nRVVZVheB9CvLOnlUFaoXORwI
UNzfauc0zhSBLF+dglDiS2vzYSerEiRASdTXhOnwJwgfHdrCd9xxpvZqielKYYM0
uGXU/8xiPROe3LRUyfsvsOCSkV0A7IZziNKDJlYC20tUmHue2WwAftEpjX8rtzgV
T0Nm4Fx6ZosT4rV/zMIU8s51rkA1iw9Xsk8AIhTWfpIwBQdSUsv8rUjgGeP0p3Md
2ZQk067A+Pbq0O9esKmmci9QXNx+HdfXSDf6uAuZisbc8jn5LVsVdOTFUDXTX6V2
lUOFaVVr/jf0TrJgKfdibeeqd9of4q7WpWo6kMek2EoJeZ8GXiEWNDp8pSRfwcwW
Nei5RyCi3o8DRUgGhhEXVD7lf2413eVkJLA3UUUvegWuwUpTKLe06jiOktCHXzVe
PsUxBrX7xXJCSBNTvcjEZYeI4Iq0PdTwpjTsrQSUzkNUPShGTc+L7zWbwmRgOJeR
sznIXQw21oBSZDCpCoJgaoRkFqek4gin2n7vAkIRKGLvoIsBN7XWs8+ZsZm0Nr4F
W/DSP83aNVu0Wk1Cf8lc8y6qq/DqaV7eGpMYInRrYmRa9cfj5m74NMftTl+tz4Ph
4GcsTYAtbR99iSfs7R0fKH7XahKDeeF/MiNZLPWnIRl/7MwVQ1reLAu9/CdSHiih
4EOEBpo9+8TsLaXT24+MXOZd6Q2wGPR0GLBtYyc7iHLgFNogE+esrxkjNVBKl2iU
SsgKlicNQKsrFgl1VSoMPDizXchWsfAAwb77hpphCdtkkA6+rGeN630W8KCbPS9v
Rc3qzzk7HFw1Ao4KNu4U5vBp9DUtafSayvYLiWc7/fGrv5GUaz+zEKCDFwbNmlq/
jFnr2jNmNhq7MjHaPdJMyds8HtEg2g4c4OnU3x1qUBjQQ0PbgUgGLJoTastJetkY
Fh5R6GhyZRhl/9uetRkPXGEjKLnh8mksvMjtUeiM2dUDkrdcGGdP5F2ny/qfUy7I
VbMnUOi8hveTM9DJevtm1avGR9wC+nXkcDS7ZLs32c3DxQnfPwBXPIi20bjDnKUG
IZvAYe4YaF3Fl6snmn2Zee9bxZMonEMriRudMvTfBftxZUmmqDWr23INeNrUqRPO
gv2ksQ7HRwigJeRtf2djyt8QGIzpHYJpAT/op6BLX5dZAyNRrnnZesU4XBBYYR2G
WYz3pUnpZa7rnA1uLLes9UacEwhxRm6zju9LUjs1Fg9YX2Hf79MikGfRkyyspDQr
q7LZaKgCiJjmQkHhSSIevrtSQtdeZjcZIys31HA8vges6HEWrSOR1o3vN51NlVx8
5misu+O5poBI8jx5Fyzze6caiMObPporyfw5LtqgSPPQFQjgBU0ESxRzJ8DXvKll
QawlbDjw2EWhiSSFicR75ffCUEP5O7DlYWpl5zGptXacEixdYg72yjl3CLm8Q2KE
MC0g22xNFnaxuVQoYCLrp5rwStvJ1uZApn+n9aGQYiyKujS3wnk/rTAQ9Qs/db1x
/itA7PaNlkpZDfCpjlRN1GFiHylTYAjgT/qzPy62VVL7UhClb849yFEoRJM17iUu
CcZDrWIl4AQgXsLu4nSBEp2VZKI5iLF72FBTqzbHIJtP4TYjHbtci3cXgv+6Wx+G
MfxtYKZuwE36v8JWeWLuykp0EctbwF0ooPTgBvAy7StUpnjZf9bEeVshblozNZxo
Ip9PtXjGBgj6sRVtQngVXpimy6xcUdC+KDtVOeFMaaDXbsGaoC0xwAXtyJ3ZPLX+
Uk3tQRQ4DqaV4LGf1TsiLRRJwjwlQ8ZoWv268Qib6UURRyn618Q2CS/8cWcAnzVU
gNa4DIAW8iB/dkEu6TwLiapVbRLyuaTOlzDap7hqU0DOQj86DP11/sN+2jCTe13+
P523uesIo/MdLEb4IFDkfM1N03b4vEGInXdWQBOXj9ilwoAV2uNDaYwHzEMIrGXi
ZKkhtFS+bYpRl1ACViAGk6zPuGwShCl5QgzvnlzUoD8IrEJIZzWMtP4K192xFaTx
QNyDj5AUbofd9d2M2hmqHhTP0DUaDDTR9QaXDwCztonDNKvWoJT+dhLqxbam4OFX
Hk2AE5Iyz7nafUhbIXXHZ61K3OIZbXg8sWROIwQiYgnX65+auSx1A3tgSkw6aVf+
HnznRjLsYzGlHQuTeR5vGx/q4D39/mFFKizk+DFUZ/62AVN7N0rPuhKWGV2lHzxx
qh5r23erbTDokbiDbyEHYFSzJaJ+1wSTxcwLESk1PRjHfiBvg8QUdjTpMh3J8Gpy
UT+AgvtmIs/z7j6tG75qDrtJa8HycmSPKgitYaEbeJLTkWrGW4NVp9NKzEc2QVsW
8xvB+uUUGnXqjEQpNrJPRlQiJJ7qE/fWT5TOC9hTLi7UYx9oQEIfsDBrJM0chxtm
9uc42NDtORl4CpC2MvO3w95B2Q7+HU8ar1WiUoZWrz6o1+r/FXJiPSq3sXWwEft4
554L/gOS+iPWYyM53Wpario+wDbaTlt/CJVQhdkAJnlzq9BSJ9kdu/CZnN2+V742
zhXoCwfn9vMoWCLejzh0PR+ctJPP+l4Jr2D+Eyqf9OgE9SnNNt4UQg8Vl97mUrOF
i2PD5Hhu+dURYOYWXFBNr9PjIqo3OncjTtQBzwfpgaYgw45hIiCkC5QxwpTun7oc
kUC9RWfrazUs6eyC76NONDRxJXrUAWHxakcLEcnwMo25WZOip/+2pl0l47AutkRC
bFdBudarfSB8uD8HBvFXQsUee7JlMZwZ2AzJGWEk+6hM02l2/WjFsr5myt+5FYkj
GzZhw+zIanwLHCxgUrgzrDUNLQ6NGBYH3SuDhO/JVRJow9hDUHR38SaoGwfKzUoV
nveLhX7KGKM38HbzuELYJ6E7FXUMQB34aU8DxV2rBlKRgs4UGDo4pBIqO3kmt0oA
JBCR1GcKEcxPanQ/7LiX/MUCVjCZOZzVXTA8LW3L0G118A+7Yc12PKKbDA2glVAh
PiJ6i0CWs2eIvm3xdHnK8f/ee5c+8fFTh9sprK6FO5Tkf33oAjeGafUIRgwpoVFw
N2a55Giul9i7Z8jJYMmwun/0SGwB+YSXBx5Aj75IcsTDoQ5bCT2CxKgMP1QchgCF
7pslOobRhKPBDuUA86xm8xHMVBaL4ie7swao69Cq4BzmRZjcNU0kUEWlSmrogCI4
nRAiMYi9+z179MfscsjzvM+BpAUdDgDehmBnTHEnh/EsYzCvp6eC1A5CUb6g3ZiJ
R9XT6ggdWf0SX/2KVmSPB4XOJ9Dx8zVqAob4S5j98WCHCefZtzkiiKYmUrAlObk4
EfS+CNnSajwxpzUMJeXNPO1uyUEWN5Q6hUuR8iAYjq//TPIkbFmlqeFSFENaLpI9
R58dzdUnRCeZoiJKCxQOQ5d5fIw7he/KXb7SAaiSbNbucjNhQwSZ1u2TdVCahrJF
Tvzn/bMV+E29KaE4DxB4I9lVV1tvn2CLTybhuGfTu5AtZGTEdgW8FVDbkp/lk1qs
ClD76ar31UdLyLvi7pcDR8Aoi7mvuwRkm0rXVTY+4Flfvi75ynMtPZgMXK2LX2Ox
ZK2PfMaW3G+C26Wzq14qQj7jvR1q64LAZjTJ8BQiR4dkgu84U4bjsi6aNLMrvUK6
oom7tf3SJBKqmSCQC/FOripRqVLPKhlg8TdxQ/7w40vqKFdTYP8I4kUYIM17JRUF
uhHDDy/8ZkNkulDTLXc6X5Ti0ydC1h7IF6DkEA6DmEKqpyGpnNQszE7CfwJeHJLy
tPYOMP1i+UVSOgzgO5ms3qRuun965E8UF4ZuXlmBaGcouodpzQsRxWUTZNDYhMaG
ztuOYUF1AdY6cXWBKuKHm8nSUfILTy3ictS0xZaP6r5Ysw4VossS8TZyNcTjuklx
tVyxnDDnIzxGiGtTwu5mWcRn5OZw2zUjeVolEzHUTMnPj3IedediGcdXP0XrG3cz
+7QqWoPCvHDrh4sQhE74SeNnBfQghAsGFRen8evUGepOd0x6qLvJ0h9U0sicCY3Y
jBwWWhbWEeNBd4BN5zrgJnvLpvWCMmJioipiGfIUkZyHXtX5aHu7tEqG5w0kzebI
5nDJ048+BXpTiZiAKx8YeT5Wt3FcMVN7Q6P8zWEuGWFtn9HAk1Iyh2fvcPSTCQ3W
E9TIhVn8xVlorK4m8Cqu09yYZCEoMmleXAa+KjE4G0hQhTH4tkMvsluooxxQ1eLE
oALU8x0T1cgSBCubweNvxzLY6qL0E1rTEcmyNv2Skc81EkG/OYxgLpOykd7UXCbW
XpnhfQ11MrX/p9zdrg7elVC7rrHWnP0H/BFIba/kdylLk62zk6tgbun6uCcLRBRb
vM0kToCprspIir225CskoqNnPN37Fb8XaDDJUdys+mX/810/8seDbBHetoOizUwt
LYMS+VLoCvUBe7bpRaPcMFlzdTlvYNXk69bNJCyg6wttk8mmQg7RDoQevYPLsMwf
Ya1FbPQUtxkfj8CcoCGyu6Dz+ix+QMp65czgo5SVGMHRbZvYbzG9sw6AnHu7WelW
PnHoWsoF4zZvmwTNGMl3RgsIyC/vfhJ+pEgfRhJD5EkXygZObr/+SNMsEPh0N6ha
0Sft1sstBqHAhpz4IOtfP/DQMGNPsjXLqnvMNMK2v3Q/TWX0VbOz60jpG9fhoC9W
snIHbx1kT1i8EdfRrrFGflb2YCTCrUznZp/gf9qMIzTdjW0R4G6A7VfFCvaNiQov
SzVqi/0toHQaoQVQE8628qv8uCHpFwKTRVIEpheextqvzMTKmera/CnPvm/dU8te
2z9xMX439u5Bx1nqcwgOX7uZ5vFzojFq0c/COzlGSLqYjFAmFl0CvDO8pYTj9bT8
JqtZ3JghrkAlzAGvGE4YTK0eA31F5XPbYP7Te/28D/v2EAG/Q6aYm8ZfebxHearl
eNGD8UARtnUn21EdfkJ7krg3AtJAxxN+YyHoEraCIpoDO/5w6S6+nCcIUtsw7AKY
xVF2VuV3LarUoq8OsgOwy42MwjdY3/tdW2u8Uwkkf6JylKd32oZJVtswDf+Zviz8
LkHHAob3L+gvGnPBbPrydn2BQDvhREjojKdx9OSSwkRVaHpH7CO8dy6sq5dDFCFi
oOAQfGhHAdbQKHD8A0Xu7bnzqKz7tEPqNvozXIvPy9yyPFe/GmRtGrNq/se7Sr0c
olfSal88mMeSfDVE63cKcZ4RMq7C3v+utU4MEnjl61MS2Zk2ZpxfRn5UmiZPSWN/
ZcMle/4JHYS/G42Fh0+1tIzshsyaLcxyi0Df5ehVcfW3isdpLfhovpq/WM9DfeL4
Ys1e5kd3xoNA8WGKLNx8tXBlIEZdUfUlWI9zvbCsO+ceySM6EDut1/Q3uOZ8JksI
vAPk3PGXFCQXOkF6LdcMphT1yJw2O09LCwXnP20VWqA3fs8+T4Ej66E9nkOChfV0
VNrvE+qo+DCuSNpqBgN4gul/mxMN7wxPvS9FZjo22bHUGeHCSerKh2+z/+bC4r0F
C0XXul5e4OnhqaMCH9qRhyEs7cqWd8ojNCEXbMdHB5G+9sLEriFiZXw0Bckkyxjd
NdpBDepM4kGtNMlxOlRwf3n5KQcsZKdMcgvgGO0wl8pzYIiLIinnbK9AchUOfxJ9
f3S47fWmEDQwpAjwY9SiR1Uy82/ZoJPagZY4/TIFggOE+9YLYcsTkKQdiH9BsM0U
CnO/VF0CNyCbMmUn7ZIADoT2b07bUdm24hrXwf3jj18aB6sgeuALiAL5oWHERyHs
eco1boNFHbYY06M47g0W6ZMl/VDLu0JlbRWQsDtkXZq7iEH2FIgKDzOsNN5fa4yj
SMC88Ku5zmntNh4iiPX1GOoeSeMdbt2MYsVYbdc+KHXQnLcagyXrC8KlLjVBQGtm
5S42jQhWHRT/FpHFsCmcn3nhFc+5wdIw6wZ/srzytf/OtrQwGJQeq9K5SGKVbOPc
uNGFQvLTz1pANHVDtweQML+MbeQSepcs8Lvy7fHHf0136nkUMjovWAz/ZJsk0BSB
s1PIW+I1B2IYY6UdrMwE+p+2J/0DP17iMjg+La0+Cz66+zCK1PfK1zmOdJ/GJ0Zc
ZUPQlNpAzMsao3Z2klLcU4FeF8hHS4dYGFC7atvsAU+w4233CG99JlYKJql5r/6d
FTp12LgA5XCgElpLH3Ha5lpO/roQRuTTjJ+LdUHjOvcWMfU1vRgdoRms13uo7wud
lMdGYzo7Z4DEnFMFK5e8rzoWHD3DmNMp3w1xG1osbFyrxWaktBwXDMRSgC3GczQG
ApqYpxnmfNlOLzNdiE5T6PLQsCd3wk8mF2VCVnt2p4uiUKVqJvAXRcT6IHdoAcE2
5Z+g7JoL7wQtFIetSJy7OgAmjkXF4KD+2V5Un4tYfQgblS/P5i+FTX1lBO6EvHcl
KAE+Jir6hXRqRQNmfbzRaPzXpoeSXTdOYQmFbhHGTceXFdrxspfMH/igy8shdyE6
NTWwc8LANkGinO4K8T8Mksok2il6azCDxKcXa75/iUpTeYD+DGmayM1yaHirLPZn
fn4BE5cOWLebiMcYpo1cj2Udndw4T3hkiP3B3bRhSGPyE5OsfbUf23Ql6uM5rY4f
n8PzenkTQDLwtjvEMqOOiF1PN/iIdJNpOO5PRCDu9fapOK3sBR5nSxK/H3WzgHGr
xGg7F57tNeHOjd8AEZaUUnmxyA4W9EnvROlqqKzj1YxqL8lcSSVdGKlSFy4XKRyB
y42HopNV5bsvuV3+wutsr+YV234jcmlQF17mkgTYJPpq3v2TweeVam6JI3tjpOMA
D5ibQsQz9vWW8p5h2sQaY7Ts8rAFZ7Wc8xNkIG8dEJidEsNaFZhaPnRxO5Ku7g0g
JAFARfY04XzBdinOmvHMkR40kiqRidCI1gOhhWErh9hH8Gdp39qfKFYJzOKL5YFw
hdCEygrP15WBwTDrK3AGKR5xDFjgIeRVOmH0kr3MQIsDqsr/qh3iT8/5Zsah8FVa
9q0r/lRSeJ3KH9HbtV1pb+Mm6yKthwDqUmPrZwkj3ESUW1tii88NjbPROu265MDr
dYNg67XPQj7meS3GSeZUs4LCpYGTBeT5LkVVqQtN5aI5JqzUbBGxCjS0FKoPtb/U
PDTi70rwTFRcVKm77I5Ih/BUWzW202c9fGKIpGS6H0KpNgyC207LmzFicomoBFi9
axi54NKUcP9sXmMBGGtXIpd7j9VtoG4R/LmkdBP9uXpUOLdeofkAJ2pmzFoyzhb8
83BO4CTmj3OyUZ5RLdwORta0xTL/fettmgxJuokGp8rSrJrud4rXq0lgziGq5L1D
Y7/iwq/1uxctBx0UZ42yXifzP4AuqviVCNmYxBAWDrcLfJaaDf1zv6xhyZbaiK2T
ZdD2e5zeklYWINeTuklqdB0d7BKoEQVoe+Kz+BG0Etukhyxaw+TIwldT3jfGOn+s
XPtf4dNe9zrF4OvjOTebej2RLxet703QAN8Rs9h5TK9LhGUqHMDlNE8q8a382kLO
GQnfOCM0X2BiyEsQli6gCrS3vwGSl6CUsL0AVw4xb7Uye75sXkng00FYqVcNVIyK
b5HHnUdySh+6X4fgK3XsDopWfla1XTXZJmhMg3QVcEmzhWOfMk3Pz+26ziAwIuOl
l9PQpCCP5ztJI3l7RBTgoQpv0yJsIlK4f0Gn7vJyC4uSRc8aUMcGhbd5+U4LGjkl
6QdlxW3VFs2SH7df5hP/kGbQH0gcqdaJmM2EUKlHt87v//wgxgYGcJ7nePVU8bPq
5CLeauTQzLBLdF+CpNJQ4FLKAQVwYcSeeztKActuhNI2kiZPx1mjQwPMyLiwhuLJ
PVFJP0pJKB8AAcPFWEtbVIcjBFtN6e2CTMIjlhIQYOlF9n2dQeS1nfCstoIBDbjw
mNwliLqWkZYXissN9vtLnINkxc4HHE+2r9jywUUVf4dSzRfxaZbgRGuSV45DeYbc
Zs4Ft30SUrhUeh8kReocTh6LpVlnfNEo9768FH1Oy/FrFQIYVWkyRwNzCZJ/Oj/z
6Oa0lIttnHGQV2bPUpXLfvt2f/laNmjh7lpG8V6VyUgHIhm/bEnVURdVCqZlQNj8
d8HcTDlVaJRYxkX95qp8c5ulrj+hNd2K03LoiAqiHuXOpaEQGbl3qMEo+T4yirvn
1wBYoXQQHpgrZG83yA6QFSUaxuXvvTTENkMb/0DTVzWca8FNyFkntn1C8VhxLMjr
hdmDtFpIsi5IvHNJBNr/LqynCWMylei14tuhnZOhPslZcV4NhGiOfB+q6RXgG9Ir
awQteBmMiDgj5G+LyLDVAHYcLo6HyYXx0M3CVkclfaB/RjvCVQ3HeqJ2HqLmkJKW
gxWx2bsE+2jzU3ya1n7tOkzww7rSqoY68mmjc/Fvu7XM9qumHVhdMqaOiY55i9Hg
taseh6pl0ADzWaYcYirt+9TETrbnrf9vIQwO+Y6/NPfRfDEVI1uhVWsjoGKWpOtf
+D0S/2+IaxmnlvyzVwoOY6whYywvy5OfYhW9bqQezS/aaM+qltbQkAAoaiKyy2BW
7o0s65AJYhjnszUKNN/7D+Pl3UfJW4wiqTxpNUvOsKFtCoWqqu0yrNVaDVFjWa8J
4roOh27/Vhhz0BzIm9K2fpsqKCoF8XgLRjXtPAaGP460x/1P3GOPKFU0j7qdQHvQ
sz4+Px2L7/GcmkB0n2pbuPtDhMI4saGEqe1SJyZWs048Kq9ZzyC51qkGAxSgCSHa
yVT5T/88ACmmgRWog0As6s2BbyI3l8HyvVGAJ5BjBO82WL/arAwLArA4fijduiCs
eZcETllshu0YPEyT6vyxywmcjHpWcxL6nvN9xBvxIOQigBiuC9Z+s297Qlpkg/uY
P4ij9cHI1lDc/l3kGuj9/jUonRQMXIcCX5WdokQpy7Xz9dEa9H2FhveuSV6mLbWF
ReUCcn/O80Naldlf9uXFiUiE48NwCNGknM2p5aqkZ401jOsZsRnJsBPuBebAJS7c
PmvviEh9U7f3KrW932WKjr4nwHEFjjoNEzJn4+GohJvlKDT+j3LU7rOySZlVYepV
9xEbCfNXed2I4hX8iWEuIY7RxsP/0ADkJmIGWvV5+qYRjXYGGyANDoa8qCLofUzd
mupwFocfGF6xiLiYp3QZWXrO3aJN8xZaHwL3vB9GUWm7SsTjUB6eymutXVQC5Sln
Kfg7HKVlF00qrWIDEsKoXnP68R/gzVRQyZsAqNHaJFCxjXVHIXO7Noxpa3uLTD5B
E9OSLFthbQeL14sHf0QwJEVfMhKOWch6ngRFDJYBZ7fJ4zL4mwD4M3qXQk8DYL6G
6Fl32G1OhdUR+z2fthQtIJXa9wL6cB2+fIiKF1g5EjTmopyJOfPUPNd9bB9zASvC
7IFQnCN1q0bmKG78gUsMtQb5wAgUcOjYqc+5tMuUmnMBCdaO4EmtgQRk7i5bTCtL
jc6XsOcwc7maqkULlyDNokvaISisObkoRttCw+vrCz9HbD9nIhQqEsoKEduF5fSn
12ghja3BToJMUahs8z3R1MmY+uMVKbRn8gA4awG2UMqCHods4+v582UkLcbt3Cbg
wQ4Smh2gQzINf54EAzqKN4ulgK2Cu4qsmYKnvQERA5QbJb4XwhQeQtzaRp4GhPp9
8uyyW7wOUBDktTkbIh0BPTB1Ppkmcbj9XThhuQcXfNV0VLa1QHDSDk/86Q8+aBKT
BmIvexylpI4jtelNBmPXgUGwKRziELwbqnIA23YFGf2/4NnXL5Dm04TkAE0AZmFT
j1822hcUbK9XsZPjysH0o9imKmkPKplu9K1cPb3FrHgUkLznrW8qtFtHtaInxmNv
62lGSbfYikTG1Ys7DhiRzXABMmHlnejO0NhCHZl6F+0ahfpMmrYWypDPAMQXZem3
WiCFCxN43s5jqRXH+Pe03BTKpbNbu+OsWOy4usHFK9EHkF1utp8PAbdr0CX0MBRX
lUxWnjKD68mTlg3+PQLWoHexKt6rXCBeYHbBaTxJ9+26fEaFDup1teFG2UwkwU3l
4Cskn4UjD7wo+vpVoMiOTIk+bYJqsvYlwkmVlgjNGbl9+xfpDYPSNURrL5hgzQPK
W6FEDlYZavtJNq8TKAaWLBhdCLyoBLiC8GTi4TgOQ1Yq6DfrZL7ZHLG19h9Kx2T4
FNDasrj1M+kWKxH/dl2UXQ49ACTkb1BpeCkaVCjxuO+FMVUErMoPbc+Z2v95DvvX
YUvEyEA4rFHS0XpX37qd/hp1QkAPcNtsWfsFO0P2cEuzg8VaUbN8x6FZuAoFrBJ4
hxr1XqyleYFG05BlrYvNpM3EdWz4AkvHOAjHszSs1uisdn9PDvWmyH0i05LeE6LH
mFMoLnL+jZsIIbVZfBxlGAOKlm6FjHVjIrk21oRIFAyohjInLaLvTv/F6uri/FQA
QQzIp7i3zbvZVudif/QCpZ08nkQCr28XsQh/JdR3QDG2eIZ9tISfqd9D6IVrdoE1
4Rkt9oaIPOxq53kxiv9EfJHQAQhhr7YL5yZ8awEasiFjTFdXs1fap4Lis11OKycd
il1COHOFtHPBG/ssVa5ZVt2rMIlJYAbpr6eUsZ7hVoDWhzJKrE8+jDx4Xs7/azuO
Fi+TxwlZ8RS/eF/PP70vK75PVB+/ci5/ki2a0OVeB7bUy+/2tjDRgWrn2Gg0jYWE
zyNzYweSbGYRJFamLiRP63x1KtsQxmRdy7G16QEXGJy5ykRMpsxNuF1rWbeASQZB
Ppuj2+UTpMrRknplU37itLpjFCk/nTmP6lZmYLPYv5mtBNIEPQAy4e31xJ1E5H2P
nQ/o/E+B04YjqdFiOoDX5YrQ2qQZYpYhAEnPo0WrTeGflKNzz7FcY9ZgbxANR+mh
HECw8HEA+yGX8cAWkKvpaO6FmPVeWG5nf8gH7vhkn007q0eeNwmkVnGOtn75S4JA
H6TDqMrHEOB84iEQd91dioINWvEdlWaFkxOrCt5X3sJAunnXucl4yeRfIiwjiq41
Kb60RYK30djiDLaNS0BCN+J9CBZ5AB+FvH3dCUMp1qlGw7GQNmdiFIjVJbuxNvvB
Vz6iOU6v2DrSgQa+G5Z+xn22ySIWSOQa1wXJpGHqPzAr8ddemlB5srajuqk+vaVp
tEI49GfHbIVbQkdtIhavc8wyYw0PHP5aD6uZk2dKE7mWI7/2qKBksjO1xOzkPAuE
34zuCeKtLDlNT0LPGb6ShECktb7ZlFBWhnux2ol2BpVfjNu6Px+k9shhKOnY8XXM
1kKU4fAEKR+rsK7LbKBY4VDhufGl5ZpG+ZNFqA4Q3cIfWJjPsm4OlQNo9cd4mWY/
ib9SARpWmu2TGX0qVKmpzb4kq5dHdogSav4T+PSHXrJNVxRGlwx1VivhA9RGXm3S
CKJdNIiTM11TU0OKCBh+F9xmmaHMt1UJSqla/81kpmbeYdDeYAH64nLiBS9JJwly
75/JPg6OfsdM8sxravA8e4FwA2YF2eKzwiGdxZaavcsIfczlkOXFwjfqZa7LnzU6
MOwYptgekEhW0DnVI7Uv3PAQjPtPbl6W43R0O3KNbo8vEZbvKVQ9wTOPGEgZSeIk
dP2PUoIc7Hs3Rw5K/HZqZ15RV+EziW2ghjgM0/S8Fj+UrZdbQ1qBpQ1AA1nCKnUD
uPcUzG0l0qVMIIlX7AH9p+kQTSkxmWbLLVtroP9F+8ymVcJ63Kkf8KqKVZZWa2Fg
dJIol04OJCxyc0xD4ug9+9TX4IrgasgYCefk3ZsrwGWFQA2tEiWatWjmTs2tqdMT
kHtnp1LQn+l3JwKdgfzleXF/dcRZUBwc999/RpG0LrwBvfWrFbOXfZPvfSM+Y6wy
FmjRIKDl4TRL8q3Hq9cJSa7orUrjT9pmXhhnowbrnWGl0yA6mXzygjUFPSPOUs3/
UfSE/DLmDWn9qh7alghderle6aUwgY8LlCADi/AWgTYN+8Gl7kC9fx/Etm70IZPf
bGZ3Ubw8ZRTR/Aay/7xPwMGoIi687jVTPwBRRY9XLXHdfflo8Kma8AfdPAhTLXKw
qzEulwWw/nP4V615GtPVMBmiGiLBtdflBvjT3k5WakCUB39PRH5R3y4DaeQ6d3xG
IcFOCIqJHTodfwOZXXPZCH/lpEANnYtBwsFOCBEl6dxCaTN0Q5d/L8E7FKt4TVO3
1Aa0A9S5uZYqTOj07iK7Gg+bLQU9oCp9Cy/iCv5UuS3grwCUWU1Ui6lv9GlhiCm5
F844Whoa7iW1oB2dxWSBN1240JWqTzVagvv22PkZ/6Qbi9g7jSzgFsZafooV8qOH
YQ7+0hcqhrkxm+ADmZviAasY0gO1e2dazN81tZ2o43/bpeNA4ZaEQ5zPwDb/TsCy
hA3hCIR6mbbxfXu8S1hPPtemPahzlDvAtFltyWRtigrbWUxb2lSk0Gy3Fi/3mhRa
MnRh26PuJeXcAWA3vvAr+y6aTQhYE7X6geh4RHn4YR1nMnEXh5D6lXy02ECjgXbL
udR3QGGByZfKOjD4PhJbzfsxVdLFHhhNLXTfgnX26mK9Gmk0L8GPNCX1cgFcIDSS
TqBuRhrowom/tSj1xIrjP2pCORe9cZxHSUsgvtkUyxlJF82szA/qHnMKPYYwWGdc
xxXJeCurHx/mehgQViXu+AVN5vnyojZLwKGdFBuLhR9rcWwVbUwTg16dyjCcMb+T
ihvP16g/xox/sLeXGnulbmSyyiNgxnZiA4OHRVvUQE3JgWKb+JniYIF8nj4F0FNJ
s6Xvk4Xi8RotQzZLm+F5UNHzFy6h9KUPKYCRugj+tJ+fSMaYpudNk6IMKcukni4f
TegJQ+oqzsQuDVUl5/gSUU5bTNdaLYDJ4zVtZv7gZH12+DCaGajL31zHUoxoB+Pw
wtgvohdzyjPuiLi9fvFO2TdisHQGrCDDzyjolk90/PoFC1QngOK1yrWWkc0rYwm3
289EAD/XPtliABhURuD8+LbKIXUx0ZlPP8SxOUBszhc/riGjm2i7YwGdECfZ6i2a
1grWQekvu+Gs1AXyPvII+0rCO3XPYmv9y21SGJKAmXy4ayH3JslnFp+G53XBo9TO
Kizp0ePfjSawYGeQ3et97el1/MRpC1PahSEgv3ZZLcfK9R3GuyNUyVoZ7zt6lddc
4PBckrS/8Rj8Ec02iGsM6Uz4XEpuRF1SpuatOkFunEHOapAN9B1Ym4Ixa75GjWBk
sNsHAPPKR4Tx9so70HklBTZEZHy0T5G4qRBH360MhFnikE7OWGfdjJWflyp2nCX/
Q6jHJGT5Fnt7OwaS8jPq64k4GUHTMlyaMc9eoej4jPxihUD+LvAdeNtbXvFpooZr
GzI7pqnbsDedQ2KGp+rl/IUhcb5juQEsOq9gUj7j8Tq+pXSACo6jPROwKenBTVMi
nxGPRvv9vttlV9/+z0lTtZYHKi0+NW8fFm6KKzgSUKEuUkwpxwn2SEnBX82L2P2p
qS1NNAWi5vHMYOdnWxYeabcSVp7zf+qbDyfNLidEeyNr50RDMWFlkzZ0zBqE0Nec
67JtUbCODtXLkYHRuJ8GvUA+FLiVnepjkl0B703KPgwPH1v8sxqk4NfWJvMpHlyy
OFIJgtoHD+JeiTDudTPsO+0OSGUALr+xCg9GZJxGP0ZMBYwIza3Z5RPYe+QUk2Fz
Rfi4xabkzVOAqHmoUrGFrb+1Mm4zjMWjShez5uIFLokN3vfk3ClxyUGfNfPoAhxf
2opI9PQ/i6txUBrl/XpSU7LwnBim8V4/6Ii9oOhRAWY761G4YLPkTYeZ5o4Gj7kx
mf+BgW2BhRo7vzSlXxU8QXO+iu9BMTbnNmsSdkz16mzxCCni6PGc3dIWNX7lss7b
E2K8xUOXRocx+jT4XWByGfVz4AQaVRG4BAWsIs99dQUDGs1bqHM7y6qtM0jbjeAA
AGiZPMZA0HnXxb4IRGNwxFzEgWrH3UCd54O4aUPtZjrlAKp5v2vjXGtZtsg2AslZ
qge6qGcuuTfNrlJayBKH8UoZOmJN4LFBs0FAkX14kfhXnf4KsS8XA36PD+A0y8VW
SGlCPzwiaMeKJCjC/z2aALJvlqzACjm5OCBZq62SHVavFWJ5Nk+UmM8mBHbCcIlX
q+n4V2F6f17r9pBOMGs2AtMgVE4jfa0UzrzV0Ad4GyNmcAv2SgI0d9YnSoi062m1
Ahpc56ElhhuYGThJ1UXvGaU/YKVt4Isz3tbPwGImUN98+Hb27RUjeKm9jST0X0Iv
MpjJ1y8WHH3CFhnGtrXXzHYgr2emo7UOfl6pKr5r2/F5m4JO+zICto7dlMtByH2y
0rJtvoBBOke2avw+VnmkOA54BwOmz++20sBQ8GGtTCa2CdYaS9szAu+5PDjngrtr
WWKNKqxLHjxCpb8tOHlnDp741v5i7YEjKxWD+vO4eOclWk994T+rj3pI6yfEFiGP
T7CWkLYOvJHgp9/l9ZOoUunynpDfaaM5KY0jS9WWJbK0t8phggIWSAxJQvHgyBFx
rtRfZG7pb82zezDlMFLGUxBMSzSlyAfeAdgYLuWd1+XcRVpt1h5CTZ7VEQffZcJz
DAxxUJ4unc6ZbG0tbu3s+gbCnL/TPEvVZ5EdTbthQcy0AC5KxmisOQiwVRz/YYf1
Yo4enXQnyKwhhLsFEfHVZJdZvfoi4MLNlXTRS4Ou53hGBHYSKiIlmu41/r8t6TV7
buZ4EWUxiWh4aOu/1CxtnCi5eahvBwlyYesUeXOoRqVPisvVpzD1gE2W6JnMSHpG
x+4YiSye6kwYy6xLVIf+3BZo7vF0OPCkn7Xnjj/Je0p02sNfXQQFWGO3dTXSt2Do
mB0GW4F5LSuIr+EtS00axeXkqIvXTgPBnxO5F7aD5KC7qr9n1k4c4Wu+W/FcWqhy
PunwOz0g4XiZaMt2/dKuU63muk3EuPPhRwzkbd79AmHcFpbKJQbZ2fo/1VinhCUv
HR/BivqdcFVkvWL3hiAy78afSU7CtvvD79r86g4uYaAcVagrijHA+isCqAv7zBUz
pwGEEnQjXL9lp4mn807qvyYJ38oI71HgEqSgpp5x0Ecp2tS/PFSsFZSPbPAKhw0e
T/qEeRGOaqPeqzi+3+5/Xx0Fb2WKVxYbndmbfmYr8bHlwQdTfzSOODnXKOCc1pMc
Mysymydjexa+s8P8pjtDGMc5m9kwmN9by9fhJE0m7Ru7Okm+lINfkJmZwNEGZfE+
9VSpHnA0j9Ma4pp+GdGzGOn34frIS77cLm0JEvRy7Kja7ExGYILxvYXeMalL3kJ8
V2j/haRpLrNsGhQ0gB7+w0NphVybNeRWEGhVsI+0aoBuA2cQUNLgzwx/5DTgYRTk
f6cffMC2COIMYXg4nPyS37fLW3XsKKw/vBHouigOmOna9iLiQtGfMAQrGt9IzMCm
/wumfrgI2z/SjgG3ctaF0N1Bn1d8zXbGwgvaboZTF9Mew7FhGfHCCvOkZARmJ92O
nro6W1WHmh781XLRdPUbr+nhZAYH695eJMXRIEBcxtlSarXa+7lRZgqGekSpLB7f
9AhH5xVblcWhcfxdwJi/ie/LxokU7aCmXY8XTwgc/wPj70Rmn5QQNHqyfsyZQbtN
Jeu3NP7llIkKniJag/8vEh434KDtFVU20RyAojqNf/zt+EOU3JVFpRpQIAx2oeS2
fhj7ji8Cz32xhdbuWv+mX9yEXBnFjJIwPOvOVIR3Qvtvo80WznD1t0QqeAxhLtaV
C8QIZqPvClvv7yv/bnw4/8+FDDMHugD9DGxLRj2Y6h2ciLBPYXXwo3LOSnsQ7YVA
1bAM1X7ZU7rJ4yJVmWj/yKS4tVIkBosKWTys63a9K3WHWT2Gj9BxtRt0BXm5ujpo
m8hwugDB8f6o3IDsu/RxMD3IxvKr9yaKKrrnkJ25IAfEyP46BiZp2tMlAA42Ja8r
HxvwiuROX4b1kT4+p90+k/OBEUc3e2aSDzKoTjgVxjT/Y5orBjOan4MSIy9CRgZv
3WBD0i20y3EH4/DlIJDjKfewRBzALU5R9ozyIsEvtLbSzDWsnsOp4ouC8ar0rOXZ
led7EMHFsZ5qcDffkNLXC2Y5rEr+Y1gCFl+a1XkXGTLZee/9GmzJILZfpXX0ZuQh
chCVsp4vadTQ8xkr6kXmA6rcOSx4QF57Xprl7OAiamIooRjTLIaKZjUY90Hfu4f3
7EkitQx1cmwt47L1YIXaJdELmhI8le+PYrNgc7tdGUsGdU8/mtCFtuSuj7nd5DGd
a4FRxTJo9EmCh0fcK9MFyFiIlWXxZezl6pGDRiDUUE9grHA3ycYysxn8vSKOhnBq
oi152R2D94mNWVDS9j86zcs9Xc+bnPwE1tuCtm1xdWTqVyzLOCzLASqBE3JNb0VA
R+M8ejVhQc9SygRaosdhGcflm7dl3fW6E+gc0PPhgfvqsuPQdNX0Wv1v8MvuqSyC
So6rd1oZZ7YPApPIlHbGfjzjxpfeTiJAlES/01o7UyjAsbhCir78auaHZsGbT1qz
0zEO5vOQ97RRzZIahn+P8iPrih8KW93w7AhLXZhbQWh85OHLFjnkEb/2xt7iAQuu
UB/tXbBRBQkCyg09+fMK7olbzt/4BOxmR8MLFmnEmGskxZboiyEoJyiDRh0ruSUU
F4yZKnLnUQMSvxK0H8lCrf1JnmmpV1utTltPjMz9brIBbGI5fUywr4jc3mLKFSu6
tVYwwttIQmC1CpHeksLBuATk0w3+2lY1lSzDBCqYxn1ZiUxTCANVU5E+r0FbA+uy
4iybTNFi2F4O1OSM/XAK3pKUWUoWs9JCxTfcxg0yOPp8GmnTpUbNZZSqOzDqz9HS
ojY9uapJdiHNNhnIdiL8xf53lCoFGRPzcrsOfNDgOwDEe7n7R9I6NvlTNIuJSXwZ
LL80c2MFDaphR5pYatAi0QdU+mMoLbGaFIpWbt5Ag/C3OjAmjKvuSm/Q/eatcAzr
m4jv5TUo0LCm1SKLAlO9Rm/iXzoFgpUcltC1/tm00UmJ7b3t//zQ3hTlA063w6zw
3p6Cmy599nR+LRn8DFpPsCre4kjNNK3uj0jUpLOdvYm3T+Oaz31YV/KrFQBU2FRf
1SNqZolPf/z2bpHR+9CNEtsXvpFHVm1JCHmORg5pDC2yeBitrbS7Au11Zz0WtGhk
b1I5b+2Lv0XVakp0aX25eYm/DEIH88TkcYJq4kHl5jYEN/QFzVWczezE79+jCjbW
QnNIHiux0bRttmdbHEXPYuzvsnmErr9XFU3PWoh26jhXpcj9DJJtChRcasKw11qx
heky+z5BrDFevXfpKfDRmHfwoeTvxprko3AhQ/IzpOpoHvulwhyI5vVNIDV86KIA
+t7r1vZ73oOGAaUOrmSvuCyyo2fjO0yUFLzKgeqkjlZE5YXMZBC+wxzJHaZLEiAc
Zw3Z/7+ZgDt9SUPPsT9AcHBpur/MZMm0udXR6HdnfAK9LcExgI0h01y6RHVK6wXu
AvEMDYX0fVTa6yijxzd4JaqNcepZhszQpL4kSFdlWC1Y59xmGle4RrWuIe/iwMUD
2yVZ8DT7FAhrlPfI7OfAtLQUj/c6LzVreFpkcen/Ym1xc+zShGspT+m+zGw4Rw4m
nyt/1TA7IN+uqgnfpf1JcoqmkQqCVn7hPBBxCmaxd4PozhERLD5kZz1KXq7qIahd
6sKyKQD6WVPI6cNjLAbUfxJ732fG7DAFSunMpR8lopmJhZNbaIvM20sgSf1WKPrZ
9ClBxZEGhhiPqDlwDfQKElS+hbHCGiBEJAOl6nVNgx6fZbTfo6aGdeAyB8VE1sJw
nI7ClCypU/+0OoA0kZZmpaIoMnr/i+3XcPlDeJcyDV8LMZykTDmRDX35uFeaGmHi
pnSMNsgHoY7nF10q3AqA6SaMR5/uHkDvjnbpIatYMBjcZZjMgrhwczsVJOqRSIJZ
q5K/pQLhttkJm346T42lvLsjnlqeqvSHIGyO7YNdQhBZ1z/HkI2WvWVWSbqxhfxO
EimsWF8kZG0ffnYq0E7HW9b8u+q3va4lQwEjC3IetZrSyou+RB3UswQKf5wKoqvz
4J3uVSswvZ6mJmSHqsxkDS7QqqDbNkdPxqjp5msFtmhLXgbnvYCuNLY1K8ftNBEi
w4HzHzI/iZWDm/xDMv6a8wBX0kCdM14zhbXciTQJz241CNsYtFbSAXRVlPm8FU93
ofvgLLzRhKj1cGPVN5WPA7J6V07/tl29/K3ZRE+YpJgtrJodFvnV66wq0XAWLnvc
iTek6Imktl5R0BoOq/6PL/xutjqEc7PrVl6cuVWGQrxhfKPmv1xb/5PjZuAc+YMQ
gvKEIwvcfEmhYBbo3zwPHJ72xraZikcG4qp6RxBMEbaS6rHKt7wwV7mjRYE2Urcc
EfBHxbbu3TF7IZQ1PlI5CN7XOHFPxusE9jnsTTmcaXwSmGvq4J025xLs0wfTYtX1
ahBMIrlwzcq5tqKiDISt3uDwFIG1n7iuHQVO5CebJQF9zDtMbhverMmPYxacynX6
l5YIOSe4OPix9EqkbrxOHC/EhlJFgaI6sJO6mQviwNYI/sc6pxhAJ86n6VEnFVXA
lX25AQE2oelqk2BeYhSj97KR5AeDV4NTvleabKvyPOaY5Om5qe0tBmtY+fcubNxM
F1yQStrV6meHHvLwYAZ8mys7Xc1BMvwZX2acJgrg14+bgGF2QU1EP1fWxH3pC5/T
6tRlmmQNFFbNk5XOxRlSrMyqQOzmYx5lzTD58PA/EWg4F7txCuJ12B98gTj9T1b/
Q/TSrO9lxk2pZSodRpxOUVOxjgi3TskCHi/zNI+6cJYE8V3g4k4fcyhX64MGKd77
g0sNgx630nfnn7k1JMHE9wPAGh3ryrVYldyhisTQ6MQTvLDyV4pUhfgCwrDhNk+x
jAUNdfiyr+QBJ7Db21bcziyfpWsgpffhPyHSRiyMY8LU88IGz3yAkEylT7s6yqQf
obteNoLNJg0IqOyxqYenopxwUoXCZre/M2sdd5kapbdOQ1+95cr1bkFFU79jcsJE
Sr0eheOgazh928D1Z9YVwOG2OGUflWCUWJpVgMrb0qymz38IL/Aarl+9u01vkqk5
QgPZ2LwROnt8hrjH1CDIGPrpSj0F4Y7C6b4OYH/WGWgobIa0MZRjxxm/bLlQhYHc
mWOe6zkuE14ZOav1uHr2OoYk2bY3xAaCZXmsReXIFkvMkW7TKvsTc78GQlYWftix
bpJMigA3no5V+hrC2Ui5Imn7Gt+HqFo7vYboPm26jPkKotWccE1VhTbU+yINBKob
tT+TKZcfUihrGY9SvJWU6r22+i49yqbc+/12kAS5bCNumSoehWQdM+c6Ci7XnCi+
7rta7BHxOrBQlu8inQt/j62VleQrI215bv7IpIf8TPXVmj1pm4ee/lkgGqK246ul
mBs/yLawYM8945jvh+XZ2TGJpqDAHJaUKeWedE5+yToGLIJIgNM/6OfXmvmKjO2q
hbC3XIce9EFIWT4KazDw5dtcv2WNbVGkcE4LTqpTYENDpowSPUqaqbgobyWp2/0S
yHcmU1uMoHWXG5/yW+k6nOlf3k0+aL/5Y0bmmFnGn0N/Svj6EOoqTpcWcaGiJ8n9
vR1Gy7MQoLusddP0GKTVPEPr0JShD5I+Meuhy0eO7iBBumg9MwWzH3fhD+IjebAj
7at/zUb5BDvhwenT6cCjPfY3VUlF4kCEVpKDYGyqL43PQpVGbt9qA+wSfBzF8UEc
0lp6+Je0R7PBAmZ1lygm1OTzhWSDDic8rJU8PH0OFbwIdGHAltl6KpAejqB/ln/+
QcgQZsY9zT8RvECRadivi03t28uW1X2OiLPxeNX8ohhIy5qcMyrpWQL+TY+Qn7/O
UZwvSzAX1wvHICUdPBuyXf2XkbIhpVymG5+fScns94rU8bYzwxNiSBW640eECNXW
sl0vBW0N0/Q84w2ec7uO80gT8KilNTfet1HSCIGM5/kqQcNnNLJZlHIkeIgIbF4R
IKaix8oFLA5wbh6kAKT46jWRwJ2CrlCYgBFDQ+B/sFR0LmVihGaAqrovC4We+MUK
V+pU35E1q3sVySQ1hba1JWdPPvdRyYYlCwXa3aa4uBQs+xx5GFeHdimTltl34SaD
LYancHjK1STtlRFkUVhRsdTnRdGv+6bJsTLgbAh/VXEXv3DGrfVGBm8QAwksbUYy
j92vHhO24anRGWLnv83VNP42aruxlRDACXmeBO6BTdXhUglYNWSrUFJRJZ7DZMFQ
MJOKXwyp20CkONy5oVJSyb6NBcqGQKLaGlfS3JzBxA8ktXr5qFwPYuHEHNce9+7B
L7mS4CEbmr+rDC5+UDGYThrHcTR4ZSo2FX2e4mapLaZZFsDsbFBeyLgUJHQBJcMc
W1LK04vOE966dv/WyYnYts/ZOO6wTWDHVhbYSMvmCX5yeZVApYV2tLVpaMsit+dc
dmUB8Al+FB/E/1ciTYM2xBFO5JF0hnSkseptr3++0RPvBJ31wYdzKqGx9ev7aFlq
ptARmTieaW00phGCdZy0M8CH9BPd4qJVPbEZ0jIruOvqQNZwhyDkMEz3d70+pgff
IEV2zsXD5xpyMKcG2CjiWOOITSezOma4+a+BZdu2ryUiuAm9qrg645fRHPHspCqK
yjAQBBE1ReJqrpe5a+OdmKcAn/ZiFdGj/0pFXEbKNvALrV7rN9aT+nVoGq1/pV8I
+ZYd0ZdWtzauoZvyrTV2GmkOlE8POueoZNhMq+78ufQJZDOej0F8YSWDfWREZ8b0
RozFi2mo0KL3jTVe6OBgb0I1gWCXwArf5OX7sffUzK5Ulm51d6utZAJGjTLhe5WL
uubsSdsXpjt8ppcx0Wh0XVlZcoCOMISoc4lTMJcjuOfJxpwUbVpZFVdqWjLmHRgo
hykF3/zMscqGDmHF00480i8VDenUbPYXJ1rLYmTBaoXNSXpZdY/DP5nk7OQvaxL3
/8g1xABiE23tsPXwqC9xr5alo5zVHh6/Cy/QFgFAmAUrwx+COKBL71oltIfn+wSI
Pd0UhgwkUnoVCTlw3/PKku65PDafBrCDwBO8rATluxuHWrHNmMBbuJKg/WzIiFk+
D0PhRcfFPNDZC9i6MOKXc+4kzTEuV90fSJt5z7c4ydhZp+8L5mCg4v1ph8k35Rx+
aSsfJo58Bt3Yi23pKBHyFLaVO2CLvIwoam4xqtNX5/4pVRbG2yycOZjmrpvnRqye
flBfDHxID3Zory9HedVpRZNIT/Y/yMiCzoaV6aO+YAK6SJjyu2371Lx0u0e7RUu8
MOqsgCr7QMH7HUJAgACuWT+djX0kFsWwZtzdhU5zRmmfkpEEFVgTnC5KkO4RlPKd
LVHJvEM+WZ2RcJ+mWUNbKkarziMcMv6887qsh0TKpWTd2ipWpih2WzbnXIaSeXrL
GgpJ770JOlNnkjcsVjK4gs5d9e0ISMigNH6Srf06YRtSfTLcfjdCdM/xZoxZRLVI
u9vu/iIIXSbLE3Dc5zFXgyMcEufKlLLQJoE/dpbsNQuJC9Jg0i3NKygMV3hCEQym
/+w9oH9Vyr+49URErXdGxGwwO7ecBD0BatiSiLrZeJPngRcPpHbcoqDX58pvuk9p
taJdwPuwg/ULW4PCVjAA+d9Xw41DKVUMlJk1MS8DseoNqpWpW0IvrFkTyRiowrVA
//pZWzV4i+bghRch65OAe0GVpYG62bzwp3hWXXWXZJu80sleXbVCbHmgq0DULJrk
s/gaVFHX58C65Q7lzEwZHRAiITtfwsYzDMqJxvRyPqjlMm6IqZp5cXKkeh3XvMEz
kw9GVMTkzz2tYyEAvrsLyioAzTCBhVVGmGHau0PE9Oav0ngjOA7hvWkLGANyT7/e
50mfqPoqS8LA92MPY37MLHGi7pVK0ePiESSeRvPYNpLXpGAhCcK3gezhkZZfXnVl
PmPHhkHiw7yuzIsHNs9TlrdeByF+GVzOeUtRjwf1sjNeASBAVFbk+lYaheACUuDL
bTJcaMW9oZdOijNP3Nz7hqbjLk9StHycPpAjeh8zbmVot+it4lIpub0GLVuHVOgN
Y34APJUG7QoCAr8jxbBXDVOVtBWy+L5JIG8QLdNZ6k8R4lkf90toOcYftW5vJRN1
8ERgeLF/kWe9DN7o35nKJod5oTZBjnGT9oSQ9529plx92RuWTKrlEgju6B53DF2z
jPrSZGAzDY+ycWi1pbqGSZbyXcIir2hsBtDnrcNW+9AQ53P5KoKwmyYULGskJVqD
pERVQJxIFSY/tNWM85rJnqqo2TcHZLQY3CmxNXcEx/UUplCRxfOWYoFL9CLnl7B4
kAQFckpb8oKea6F1MUP7m5FbWqwp8jnxF08Os0YiFJ8FUbhS3/fxhQ/UZFsFLOSG
G4dmFNU+cHZ+Ig9avqv+n5G7q6ejqodYcMqGndvFkWwF8a+Fn+B3PGE6eflTXHmD
eDOGtCNH6mXyJ6L9rDe3FHWBIWhmiwR0P9YR4CAVKoCONpIqh3sWTwsBrRK4tZNy
g/RFoPa8Tkcyj0bFqzZ+Upp7GpJMw3JN9SsXFHmin5EdWzVp7qtokQvSj8m/y8FJ
6d7uHM2wByn87lQFrKzmrS8hIaa81jureF8/c80I8qEHn1W+ZBhKjjgTJRK3YNcS
q/62NUpHzQv04oUtJPfcXxOqNmSf460OsmOT/qppykB3E/lKr/rVyisJmOWKMk/W
32Zz87gziSf5izg82s9wurv108k4yL16jFQBW3lXyrrrK5JJumvLbmNF7gxH5eIy
75nrnKDCE2nKjXqkB1qnuQ==
`pragma protect end_protected
