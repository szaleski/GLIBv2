// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:51 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
I3gS/4HHFZ/p2p1b70lOhYdg5zq8WcqXMIRumRf65v8sDRhngYe/Lbm0Vcz1ReDG
ZHAd/rBW8DZGoTPB6+4kXug64z4OLj0bMl2kVsIPx4Itzn1WkV9chuykJ4GMYpii
iIsWTclqM2rTNihUAGeQZQsYyS5P0m/HP0jYo3P2kXw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6864)
Gn5tdgimC+XwsYr+TPm3t27tShDr9Qujq/rXI1N8D66M3kAFvoZx7PIKMmReUI66
gPTencmf6QL5okKw4jTs29zHX3moArd+Lvk77XmoGF5KTgwKzsz5l8EPEB5KopzX
Gb9ktsIDQg2NKginv91bbk4EjEoTtMQOrlRHy3yLziV1HwT2E8ZRTwcWCCjwLrwl
u8ByaDJ3j/czYlThCMEDPBKwNsruliLg8HTpqiDzibws6DIJn5PWr4IG5YyUcZBm
dwMeqpzzfUP/nvhkOnV2oAjbviwmkN+7xuXWNalHK8ZdWFLMjyQwf4GRKMag06sq
MOlAihzl82g4JpP4UNFimkHJyb0UyT9I0mFxNy8HS51okX2OCVn44Y+rUbNdMDmX
sr1GQZ9O/aeNbG8kpfAu9F5M8aC9aXduutmEwqWsY0txbSx7cNDWb82KCG0mQwVI
A12Biz7pr/actSMKB53EvJQs7kLuucXyY9IZ1uz08mRNfzfUCZh5jWolXy2bdfJr
Y2EcjauOUt2oW0G5WTuWac07NZZqSkNzYVx2FM/Fcv/Me8vPWYgCzZwj1KNQrMG6
hbixJxpQnIqDgJEET9DOZ5li0agNL1s53a99ZY3CztL4ryeNkATz1Ru2E4szGsMs
Jz4F9i7J1oAuqqH0dz9v/PYTSJP6LTzDIXq5sC9RzR4KpsTkmtyMq4WII/IpSSsp
vkpTfHekMphC/5YTQYJO/ecdzCvqrtnIuc49cVTzyi7qFiRUN+fngeuhOoBHZRqn
Iz4BymvuvQVE6+T6GfGub9cvbAwM7uFiK2xNRuDDDddYRu/AOhRLnXl3DA9y7HfG
IOBDtvZlx03WfNj14zuiEBQh5aPp1wmXEZ94witt1gQAo6pC3tK+HZbrmlcIriby
Nq/nvRp8OYWo1v23fJNJhceg5v5nTA12BK6qVCLMGZ3j7hNFZSfdunfjDGi/Szir
zTNk0leqz/ICELAWNdPVZ8Rco6LmAfm3dIi1TE5gOSj167N1D3kBI616nAVD14Ze
KamI3Dbvbvs2Zv2kjzjtj7z0ZyE8N4Ud9KJdQoQrmyOHIz/c5iwV/8N9HE7i6dCU
j/6LyufDjHGYtxluhJLem5AgRkkpm/rF0RoHcOvDR2ZBYcuKcPJT0wTnhAafXV/E
4ZZNhFk1HdrmSZJ+yWdueBEknry3KtRBwd0yxPcdPyOBp42xqGSYFrcoCAW4N0EN
H/TUUzqL53gEuVTvMRnSCuUV6XzbDesxQvAgUF9VOJ/N9k5DvDb9mOaLEn19yvt6
NgZlZmGECETifbDuFOUyB7j2LhD0d+LpA+1Z0PqwCGNTk7BZq525hLzkkrbPrECN
zzL9Z4VDOzpig8UfKxojR6/ti1jAHzFpwvj+1XOqgZgrKJgG9BhTOAiz5CcgPD2s
qDeBUpLY7Di2KTY1J4vFs+OJIoFcghF7IN5Lg4vUpnKv+BmzcT9i/EzrG5+h3U4N
8LajVG/4tRjmz/ELKXsxN56X1IxZK0c/oO1cYrTl903+h3OvMhZj9fiNMt0ozBUG
SvCQD1WMNoG0wZqa4mVMVMmfaJ7HC+EBsAapbKoLUr7VjCaw+CigkxutNxxMx6b9
1dLFPXUZLJ13/+pw3bs3cpIXBzb7Y0XsT5xPzDXNYB+T+kgfvKwRtIofx3JhBxBi
gylcgTCoiojPQnJmKb43UE3cTnF1sqxexfqaJzJ3imqEZtbr+77Fj/3eWprI7QRJ
NLlI6ExDougN9Ao9HOsbq/LB9/2NLkIf9binr3DRQ8Z5gXZXK6Iki4XotHF3SquL
eVZhNHy6zPqbawEUv21M3M0CF28h/rpZKdRCdnhobQHJ0UeMv/rsZuyI97nwKyiu
5sVshYsK9mcyvoTC3GWlP01PBIU1AHf1f+zG+Bka2zYiJRZ5Q8qqgWM0wjRaJONN
jw0xCJlZdmZHC3WShSTXdWiE6y/EeNZMZ5qY7olyYDrGHbPqjFB0OQBTDDgrf2D5
jfpDupumHz3A3QoY670FM4K7NtggAnjq+CTqjvV82ZQZe8vlgIoDZmjcjvS52y6j
6NHvOY6HwMClxUftyq9KorxzLZZ7cqasGPupvCbk/FVgxtsEEEEVv78Xudm4A9bZ
YXEFZJNZvSo2DAL8RMRhZphdIktXiuAxa7zKFxmtgtNKWqT9uLMcSPiDATb2hOD8
MZKIAoXPyCYx5vzkPh8mnsSS7PwKvYsW6A09fAqxS56vTlv5Y94grBiAhfu98MXp
OiB47K83SAyIvhpz0Y3NRJ+01/Ns0KqDdjFYag+0Ie5/EYKGbeGPeegtdBL0Ac1n
wykqJYNhcYhyuKP/wQS9fpSof8OEA05EN/jF2MfLOYSekpNt1RawUDZ+YjtRBWJO
8dTjKYkkmdEdY+8u5lI0wU0lAmMQ08LuPV0/KPU0D5S3O1AWFqJmaaARjsnBHmif
H6IGpOUkp3YD+D+NVgWHx2qkNUGqTqlQ0eD+8e5MJXkwuHUnPH3gElMFqz74NrAe
c/BTX/fIKfMTg5EI4UZGNlMC2tAYOBtMEiso/V2FI6+A/ClbmRo+AMUuqzuV6fF8
RVEZBQeqyA0dHWBPxSOVTnvLW5DKbbBHohaPJm113ZKwRy5/1CQmnfZiu2jrawsF
Caz+8tJyMKMNdN3uCi0K8MzTf06QX2P6aIdjrIfQuKUGU2dzQISv29R1LEwJJfcm
32rQPAOIfNSCMdcsn2wxQvSf9Sw5qnxfsXOkIv11WiXixKAGx5K6Z8884QdkKMdq
M4KQinjnuO/fN16ba0f1J4TyUu4a1am5Q2s4WeX88/NitSpgO0xwamgItHY2Ggd3
Kc3+g9umkK6V5jmAhHMOLu3vGV1a9HZnbW18u6qyTC/0oPj7Y5Dw5djNdoBQaFNf
v7EBKVxtQQNAbnKazRmXefCeJJ6JHYNXQ7SBXbbZGls3otluIlsF0c056Mn+4Gvk
d22P8r3U2UmeOkxo1hiTjx9Tlj/PBFl7HG/6MJlB0jE4peB4XrdRoinKCwlp8LAd
hon6nAFMpsp5YA6Z7398AbauFIWEhl3+I+gB6pjI878UimVinOIOcq1daFbKprxB
745tQKdskby4gIp4G4ALt5jj2C+NDNmFXyh36D0ifipPPRvihzF6Y70lAuB21eHy
3MCvzWc103vmFIXQeo+/iLyuyrLzDXa7nd3g/aJ/BYVYwQnTp/72+w4NPeGUVzew
63U7IJ+74blJmec7UCFsUr3etbgTdHdvUt398pHICy8iGDATCRxY7qwJQuOIWNnT
ocED2QbueidntdDF4Uz+YPmVs1bHVLbpYVNXe5Bfrme9b4WgSZoZAkJSi7RwF0pa
3WQ8pijNlRN9cM8bjgy+csZj2lwr/pW+kVQIf4W7X5b3rrB31weu2y/eYCICDS7i
grIwu9eLPTFG6LryVMieoevirBTQ8D1Ygchj5j1GgghmCc02aLh1nktZUHBUceDe
uWdm8qV1D0qPVjKQ4Iih/eov340dh5Ai01XkIc/u2g3wT7Rkt6hceTAMOpGdOUC7
BgCBrD4QOIC1ITxglrAPp52+eFG0mXrRvchf5bPVVMSj2qccNshW6T2X4oP15NsB
tCc9zyxOPviME817vwpSI7T19fpNapjek+QXOFVKwtpDqIImpYYHdmaWp4Kz7k8c
RHS8rNBdlH7Z2JvmcYUlaGq/v7v9X6gR1dSr8JfOVAbPHuaw+auoZtLsjUGqSK/e
Mimnvjk7992t044NWvd1YRRZzfwo87FRVRlyD5tzHYkulksJD7sSye7Xj653VA3/
vS8L9B6Zt7tyrRBYYbgeYmUnTqLmqZ5VqHkf9l+I+U8EznSMDDqmlsAHFZDLJH9X
8zA91MFhim5LTzg71qakbh+NepJYGIlDlXRL/6V/bMFT7dSjAq4Vyh7uL6oPnXia
oCi6CaZsMxe9Jsc1Yra5kYNdXho4vsTU+bXPZjmW/0QLWEILQtHC1ZR3RASMMtYA
Ipw0SJuZdENh8eKOC5VZPE2nXgxMWndheEaJZ0L6ymLaFrD5IuhTSZVxFf9ItsRn
orpwhGau53dZQeYrPyiEnRFUX/sjm1puDsbcsVSemJkg6kPq/1tkFLu34jLsW/rT
xjCHbtFlWuzQpe58DmoxfPwNS0JSHf4luXx3lelUXS/cW0DQ02CGLuaGzydzUk9p
7TrQYmy4yJDiCgk+B7LbsRf6xEgjN1xLTEWQybx6P4E3G9jzESuQA73XkgdevRCj
/8ilDOuZYiJJfN7ki6Z2Teb3Ga9NmMRFytA+u89k1vE86lxUOvZ/Q92zaWzk5nVS
d22q2ALBIeU1pUkUvEQY7qP6/S+WWuqw64vi62IUNcLat1je8TQAa9yUP//hsRxt
PxkY5NpseGzuM2TzRsLDacsi2OZaX85K6KDoXiCrJuswICSfp1J9dfcjovBfHXi8
hw10zTwePwUaB8yekFvVVR40Xge8iYI0TuMx2UElMlNihsIOMaBO+PvlhozN3oPT
LIdejIsLfyd1D2p2R1EUKMl/NewxE+YyqGBqueRii/cQbtOWK42HnX2feomb4cx0
6DEIblc4x+elz648tYgeAybLdxK0FxJBQ7S6afwtKbvCJRsxajRrQLfR+OPAezte
z6MZhB9Paswjia0xwYCbFF6SMgXipJHs46VpfKcgwuhQAGy9OJwdjAa1+N/gWphg
p2LWZ5s3++ONfQ34MumJFj1Ji/UjaBrGDHarW4ADkrSIh9gFIqa5hD478piANlVk
UefJ+17q2i5kCcQhRnV68eueDKZpNvaHWemum6SqlgCuB6CAJR4Q+XeLGuYHmCiP
7CoP8XM+9B9fgyEuyKI59t8PBXIyG/S/gAABRTVIsGLl5lkAX8Z2RZNjVk7rHmlx
dgnxoNy7/+8tHHxyTaCIbwWrnQPic5FMqN1mdUEa65/4xpm0qmz4wzoD3SBz0U18
Vxk3mw91jr6lw8tjoQZkDbw/dc8rvInqjF5SijuRXzZVkBex9/hJqKDVStX2ZcDS
DFY2ZeFB1gqzRYFMYOKtK/YVUUr0sF1eUK7wmNqNtvXADkJZcn8zErmhGPAYGxfX
tiOSAxjKiUAtwKhrgZJJhCvujhYYomYXoXvBBHsBFJkGV0DoKKbCDUBRKS3Y/JBJ
Pjxjl4e5wUxE33gR9tJgj8Ges1FuwHRmJnaxYKBXevsrCje3pzDrLiap8votm7CG
ivvuVHMcd0vHkFVjFDK6JVHzLEDuCNkUxcp8VpjSwet7s6FhEdB69cOMRJY9b8/D
12ZLrgS7wjbwEaFP8LEETGQqXy47Kt9k3+151nS9JJio2mh/AeZeg87Ze4bC6qKX
D5Xv3L30J7P2DdXITrhY8W+vau7MX1n7ezaZH/aWsQaOK1QldSscn6rtTYqJZk5Y
HC4/rac0EMs1M4x78bkpT7FmoCxay/Lr+3zN7E852Xu+xPEcnEbRP/SGeuyIkB0l
punJTElEHZb4BDiEXGyqlzrG1n0q7/6ai028VFk2ZILg/yOaNNaC3+dq6cTbzL1j
CdEj9gwpaAovyCzXKA1Ibj3C2LtA04vF7akSbLvRFPzwyhqaGSNTI3D4hAZmfGOv
TTsU+86If7RQLRGlzMHX8r9hgMSY082FAdWS1NpgJeSvj2rlRguu7mPckRhy8ns1
s0TnZ6nz07mLZvA/H9hJpzCAjgty0VbCqokhbSzdy9lSNBmcT2ivAOIF/MqgtUYo
/0v8NCltLqG/BPcjjbkODgL65HoLv1z13WrgjCu4A7ROd1Poyv8y3vCrY7ppctKJ
FXEIF0cIPA3jA3y3n+PJXY7DD74rr1Coiz+/pqFNXzyviQru0AlsjLwDY5py41y+
pi+vWtuX5jNAek1BiVIexc+bgdrgzjh+gD1gQzhyYSMcTo2CR0E1ZkF8euWye+AP
H8U03TkktfI06v65OBP8BrAdAZHdjGgHuzV5Cd3Fq0uVFZRu9zDMFKvl5HBwm2WT
zhprD+x2JDf1yr2i/arWO+4EO/b7pBMZUx6YCoyF0XBn2ZDg+o6Yi/DQI9VhtbDU
vFKa3ok36UDmW6Jnc2uijTh7kIXgF9EwkN+TcxfX+4h1H6KavJqyb/Mb6m5sGYPC
26KRVonVMjlfWEXA2SeSCLhZjkQeI5OrSdh2lYtehDc2dDBV/fd9etkVBpkB7Tw/
RJg0AjsNDY61rXHhemyBaQuzo4toCMEcIt1tFuwT655hoQTGIfG0Vi/HSYKoWFOe
G3v9GJAFVeMxXDjpuB4XCYjALJAdosVr7l2fPs6EHoxjpAzyB801iGQ/IAdDegeM
ynD9ug6wSF59RmZduLf3EB2JTKEDaoOKyRngvOUmN6F575wN0+A8yE9TmITAKDiA
w0oNx131V/q4hkgpodQqGw7lT3eKR2vvKZ8IURGF+gNb0lpNYv73k9O0U2eAUh2m
YpjreGBp+MxyGPS/PV/yb/puTK8meSlbR2nfsNlvwsH7DU2zCAuuBpo+JfVNTb4f
YEmH38zIOlkIYzP5O/1BACibagFYT6HA5q+dBM8LgkoDaRya+cTflqJiLyAb+YUT
A+aduUctbgxyIdtVH8Xln1hrwWmJDzTaTsApxAGX2OZ9vt6pDoCJf5N8mt0XEX44
csHW04PYxxok0NTEcwMLdrmSYogv7LUB7m6Wvy1tyQYBFbs0F1QN0jX9lopS+Lxd
L8zFX1836CcDxvwXLU4+luGKB7J0PXLwiOANa20nMc2Ci6EtOkZwnZvqEGREcb5C
DdF4/9jgbUKJYaNjHl8btr4AUaxGqvilT4WMY8AD+G9AvQPsTd4zno2K20kWA1BM
LR/96TTiGraXP2uqukbci7ZuzIrq8uN2d0mlpe37LaXzioJIAihbSQXix5/z5DNK
2yYp+8voXKoUBwpOaLWAKGkmQZQ444ElEfp1XKlJqXovOhT+gZnJ0a71ZU8kmQDa
sMYCKGyQOYKXG7zkWnR1it5LQPgboCMYJ0VGRwJVctqniFDuI9NMWL4tw9d3Uqzr
kU1ZUlTztiYHiDWZbhRCLIxx84O2duMtE0MgWp4nd/IggmrFefQfZUktNEy2NU3y
xn8n0ndFdFMcHrCX25FD5vHLSGG2MoyB2o2SbgQVfsY2lbr+YQpd19PZy2uxtZD9
Jva29NojUiVKEfK9sw6gvC+Uh5qXJIQYGu28wMCrJb0sWNHLKheSdGC+pvwylDwX
oPe1B96LlUTT9v3+oYkopaPtOQeVvgd9jqGnxzq5IFJMlKtfKXaET4ddLzWG2weT
SbZ9kklndVjyzOigoe2w+u4AGGFzXuSWbpi9VgZRs9ZKCazNNHubpzdlO1xoNsK+
tg1RwhFcfxyn0do4cRl9PTHfUowFs5nJ+8BAJBvP6FJkSWhEJkyvsNB7UsWx9cT9
tUF6iKYLQwqt4/z/5En8iVUpjg2M0RiofLRb+P6iI79B1E+yx32/vy90B/RcYo2l
NcwonBzr/R43SbdGTzAVM+2kF22rHLsr9A8gRLTA/te6WrBjQ53d9os0dEhL5IOf
wPFzYy0zUDdVvnCwsm3wsXiGiQ7PZaKrAnxagE5r5GxPPrz9SvsyhR9okKQz3ATP
2Tm92FfoIdlC2jrWGIIYQXzH2jbi642p4BcvlWcLDHWBBN3wVZh8Ol6mtnphrJlD
C/K4/gbIVuYum7NRwuR9Vev8qSq1fySTzx/xvFmiR0eWTER22qC/q7XHH6w0qRPs
tJs66KOEm2ZseC1oiTkbyj196Yc77Sq6/AyW6D0x0D67yUdn2LYofDZlVKAo/jt/
t/in39rno8m1LPqaDx+WS7zQE1sOrKJNTRmvNer1TJodeR1GeSxyUjB6OvgCnG7I
5du/fekHZkyYVHS5F0oJa7q6o0fojJHJ97fmwi+DfEhzqd8caoI304vW8+VdY7Pm
mprJtax6XTRAzb/oGJDSTJvba1Gb1BPfsTlvV04VU9peAbcyEWZU6ok1ze+Ned4h
p2ehzv9jcKgbl3+uZGmLJxdfNB6WJHCSQQnP6jDpw2lKqNrNIr2QLRX+/PimzVGj
cAWG1oIJFmKkn/EUE0l3jWaKg+NRZUuBp/XLQ531mNO8syhHIyeXwI+zDbhn7SBW
BgYFDgWK/MT9Gi++H+b6ETccq5ecOjNnf+cnAHwY+JUvSZZ9oXujUIJz0CCQTvtc
kirOQAgf1fwRAOHtrKL8i40gxcOvC13E4g5B11IVx3XpdSOYnLv32AF5DeyrnccS
OBggB6PAKoJcKl4J7h+5g1l+LqJG8m7mWvFIo4k/WrYZKYnfG0ZYGPoIzFJoVPkp
IV0ju2RQjwzZx+jCZ/ePw66pg4InSiITC5/6RAD+UwV9JLC2Skja0I3dp27eh4w7
pSSOzFl//BtjJUAUhdDcGZnkmpjtcoFgkF9EgcJQt75amI9jllEHisn8J3wBA+qn
Pz8MOx5hQw/D2kodySi+t6ZWH9P3lRT2GEqXaEYxz2zbPHu+ae/2FDttcz9bJ5G7
LQDSmRqImxkrejETt6g3EOxg0zORMyIPizHdKaWNOfDJpt+01md2ef8R3iAhD9PL
dlV97e8XRSoB2Le4Qp44GAD8f6Ui9Wjcsq5n51kX0PwSSGznznA7jE+ZozOOY4LE
+c5PBM9nh6oo1X/dAGQhfK5ZDIFPh7PFOXAXGS7s+bGhB2xY8TOykbkTj5x1zACF
O/pFUQ0e8Y+BX0vKRsbZCeUDl61i4/TPVQXbWqLAkZlKXfQQDl9pIJMeN/RuG/eL
RKweVeUsThtqCMFlbS4xZ3w8tcAU+MKtEEDAl9JiiQbwzt+j2irtdyXUKkwv8FAx
/FnEmqdRmgIYNoPR0LCowyjvD0q9dxsDM4KRZa7Bry+3QuGCkMP/N482k67MPhkL
0ha5fsJ/UKIRfRk0wSMzE9k5hPCcDOquhObeC1mbKrlN1nNumfy1bLCnmTZ6MCcu
6O/nDyhKaCSG853H3ErHeg6xtGkOK9YyuSk9fivPBEn8gD1RlWJZaXBOTlr+5sBg
FnVZwqKMVMmzdYnGpMJylJXUaCdOCiVGemSnn8m+IQEgnMHUX0dD3Elaak7RIQU9
bfEfcdMx7lIWB+ffXDU9o4GJl4m3y43RoQ6wmMisvJifSmSerDIbT37mBX7xRnbT
oubsea7aHeuMkZZbpg/Lt5EkDEvWcA8/mZ2mzh3mrPfooXxYN7xHwqTsVjg4jxF5
`pragma protect end_protected
