// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:58 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
MBAg7hJHHz2/qO3GWaZ5I6Svsu+8fOd/herI8Fb6BZkF8tQ9YWnNEsibqv2g44Ul
b/vdVlN23TdOieJwihetGz3txJP65IUKSA/lB4nvaqTmkJ2/IppypqlDMofJ8ZBX
EfdPhKkOi8iTsBokHQ3to6pKjzmOJ2VOJ5kB/5r5s2I=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8688)
0hGc0x2FJewyG1fagaTl3XaD3AgIdrlSNMTJ0b7mCDRKcDU6ACUteto7WJG8K0SL
OGsZc9vREZlIbInmoKwzjnqUTGYVumk7U5rpdF18w1slwEy1GQN5cHxvAL43MWLH
ksjOri7IKPUA0remqGWF1lyZ46DjxCGycgDQ8goQ9aFlMLfgi6gkvjIPz/1zoGIW
eep60Yp1Ey+ihIFxejb+HRJrv4a0wBTspLDUwEnHxv6P790IiDYT/L/Olnf7bjx4
oKFBkSjX5AW/MbKVhoOynV4JUiGixBDPKzV/prqyvoRvPLqWwpaoj6gqzoqw/zzQ
EByiHi6GG2uzkCpZ6/AogGwXuHDXUrU0g/aoQ8SSmzRLrqQSom23YY+gz8fyutCA
ajezSQk8WSn8bmkRxePTbLFCnsAzdieGaOEYEj0JKsu7HZy0GITw9JydT+tJkK8I
VgHwr3ucjWs8azYh/22Gjxz8V8RrXIP1sXsJXcaX42C6qvOOPYz2xQ4vHYm2DwPX
HpfSOfnANw0HcivGtz3tD0SligrqTFCTUVLQYuGKoI8gbt/30TVu4v19z9ZpF48K
Swi45B1F6lCWLmu9z3lXxH0cZ7r8qGjwZa2cHLG+kK7MoTTQajsGoXrrKsnzYwVg
oL9MeONkodD0f+9ckL9l/m4peQm5kh6dVm88Mu7DfS11DhxAk5KuRyVgH/6s53QG
Nk7IR45XjjBSowwl77W9jmdf/jc5QnoOiBwaFldvLVWpSSi7xYK3cMOkaZJlEeSu
mrdukUoqadIG71h+RvMIO3glnzIbSGC3+yxtpoGcsS1Ai/Fw4tlsKClp68xTBloj
mQOkHmgQzbG3NEym4upkiz5Uz2RPpAsDa1wOaeA0MYpDQHeuEzs6/x/NL722oB1Y
aKD3buZabl9S/BxNtnvBqc4dGVKdaHOMrk2mw9L2tvK6Re0S4eTn4S5+qf3X7vf3
UzWLTmhwzKEalBnrngysrW99vYEXSV3iYueIEDs0V6tqOixU94h/Jsie+70dvnpH
/fpglXD1mdtYCHmM1qYGywBeJHZnqbqDEqR6H/zgQYStkTdQTV7cymc62nsEelE7
J9yl7hyjeTqUngU6nzPcOjDDkg2qghgkU8Hx0pJyp6Aub0YcUnyxijPlhRbWU0+B
PGfij06cGDbN/ceinpEHUhn+AiWg1nrWuosQ779/Zk4famvvjvSx36MUtA1KGrBK
CkYMrCa8xAFlrZd7w9v44HgxN4gxBMTHgQAaWfvCXGIIO16+oCTo2j8Ig9dtFACl
BViCAwjZmoRP4wjZ55znYqyLFl6vUc4gssCMQIrFds2SKMKaMghqoMuvpitcYqFO
Izqj+tBzc1fvx/8pMZctvo2Cr2FvTiNQ7W22BFQhfq9+0gYlJApILFuVPMfOKC7b
MFhDvo+PabnKxvjpJN+xMyAY3G5wgwb/nRGReXgUqkQI6zVJeyIMDY4knZT0Vi7f
GrLY0IxloR78m7MaDvzuLd4/4oo/jGSzad66RpEE/3DCFG8mPsBEnh34b188eCe3
z4O3zYEYwrHYBxBiZl6zLt0BogDrnVt/Z3XhDdmi5J3PoMuC+eq150L4/60a5+5B
onJitQVoOz55uifOlYnKLPuPn90ErY9KPHgHkyL8h0y/lN/dtqZHZMnUZ9sSiucL
bmZchXTaWCdIXiAdIiXzAFYShLRyuA4L/YtVTJuPa0M/+/zL73dSpwpa3L3QGoNp
/PoHmJ0cFFbd06i7qQhf8CBNNUndBBKNhRiI/k+kYVgB0N29dcfOmXfy1ZibBnz9
B/+cYIeElJThzD54ZznIDlQwfj9O3aaJWEdF9+snYXuMbRIYZv1d0bvljJNnXKA6
ahEDYlH+dx9bGq4Ari7zh0EGtMiHVSeAAGOnqzgCOjnHi9wOZ9SPY0D87+jbnxV4
5+ZsPx8jRnY019BKoLs16oJDGFyVxvcht5kEOCznryea64dWcWgZ7YnklY1Ebmas
ynNuC6zEcPK477XFKYhJfkeJV9nYpD2uJBmNHH1t9XsBqmH/3IM0dNuyB5DKll7c
jTMsHeUSmPKIGoDREet+irW6LK9eqajCTpunOtobpHOnxOx3FlMvkWkcptottNzN
3tZBGS+GqdL+07WyWdx9Grtr4vlW/NdhOUNVNU9jB/WVgTQJFrftvpUlzu7kWNqZ
s3sriRLgNrJXA/V//PEd/E6C6MW81oHo4GbaY+EaUZC4vXoiUtK2jf75X6H1tkRm
jn2X5usNLXi5aMd5GnkQW31kOfCc4SUOzp1KZMlhiUtIzHdUEub0kQ+kei4e6lbi
EtZs8dRaV7htwC8z4rgW4Cv1onv0HoGQTKnYu+nKomXoQ89UbR01e8gjU9TgICtU
Uhd9lQ3cmC0Hq0jsF+R0HJHpQ48tDtKuM3OR8LyW/oqsMEoRqHs/XL0BLtzjj7EB
D/G3ob6zxEfdN6e9/2J3VH26oSQlmMNGaG/Sca7X+FOCdJPQC3zCvr5d6jn3siQo
Q+09kKBPs9oKOl2GQthLGSxVxvb9Ftd2NrGNfgiimPFDoFAYRkm1sCHZIyPTEkzN
AeaUuv43L4qexajDH0UKydjIMuVO9/tPe4E2KYS6kuMnzAyGyZjYPAJA+336DKpO
pNm04vHZNf/NyLQVKkt1XDlGAZ4SsKZ36kBMLEF39sxFocbQjNHxduefUaaLVtTR
DhBA1YKQP3gXlp8XceW/CcbxRaUEfI2ViGR9/yTzv+3mcTCrOVwNszNfFj4KDIGX
xRBJRj9SuOn9TMK2pJwWbSAkk/3nRi2zMjgNXuGy8MufqyqdOv1WgMRvsdM1xUNF
0vcLafIIPu6V5OwlbRwlpLfDOExLh5IRMmOqLU/WslI5TRu3v4Vi3RR4wRCJNGwE
bHW0fsj6nDD758MGWOjrZLLtnq2QNlvbikeCOwjBTBquB3b6zgFE4Ik6xTb7+MJK
sCHpr63xHH0Y0ToAhsoML4cd73xUCtIYSjYZoQiq8tyfPJs1V2Fm0XN6p9iNY9Ry
HO/X2B6UyIIayGd03HsyBCQ5mjMHo7w7l6d9+dwKH+Y/vdOWX/lnV5JzKAYiCOTQ
COre5xBq8+wngnIdqbkM6FC9NTpBIDYxkBTfYqBAGxZA3E4N5DROMjRJsh0Fn850
cBaHFgbS5PLdLdRjkpaLGY5fpxT7tSUohN7pW7RMcOER09Pkrfd3NAfqZJPUcZtQ
Pppdgj7m+GJbRTFwG+FO05EKyAAJwaYMhfbaw2z5CP1MR8GoDp9ksDkqNPsLY1f5
IX4hE7zSi90lFxpAIWkA59P3oA2no9wEy0VSiLE6AC5Lc7Q/Iad1hTEyLk2jiGg9
uTfl9DnVNw5U+qHmAq6kXoXHixI8RHjmw6A44W5Xiy9eLBxZuahM4xG8C5IkWyQ5
jYRHJ68mw8jtWdb1Q9BgoZYIVu/Y8Xi9ed198x+51ECaY5slK5CwMBgDAe7uqgW0
qUgTBeyW9UF46d5pe3JwiZCqW4muJ1iw2fFp5opcMYrKHsNUbKYFslIZHxViROlW
+/oSYPq1ws7hTbPhaVmRlNtPCM1uV1sLW/WaVZyhIKJhfI+LqQLrZ+/Gbw4p7Ql1
iu6vyq4bblQ9tgqDOpL6gxXWs2E+dYjaNjhW/XTxGMKmMWhaY/5nl3LbCZ24dIDQ
P2X2Gdfh8vKiZMzLGgCHO7t6oy/3Sk0mw/JMQuSEoEBDQ6Ut9EYIfMLLVcSgqwJ2
Tpai3DVq478L8LeelUj8J+GBu1QlLdFn9SdwxjaUnJF1n+qPwPMlDboxCb/C8E2G
jmjpEDUD/v7+vblL18T1GMrqilDTNCrpzj11jw7HKmu2IqkdbQ7krUMlA7fOAe1N
0JYAltN12rvcPoDEco5XzMWCJrNkY+Rtie7YOq/suKtPkh+GJ4LDg2ZhEmKFlA5X
wBh070RzLLl1J9LkFT7RFQ4UBUq9gm3VD64vKKnQp6xK4sHjOwgSmpCyvDZE0NfO
Z84Qnuzk2TaYyhOfdNSFt4LS3DzlVhNXh+ARxuGAjvWjigAt8Ow1thrqraEZEI3Q
ugI658lAU+PGTnTihzcXgN5QDQDvoOEksohQZWNmH+5UTJF3qhB9nK33Qzvzm4K+
jhkxREOrGeKpssDlp3kOi0gjZeIuKgL3o+PYvxDbwt/M5FZleMD7mwLd3FoXUUNq
2ubPciaPaVCBr/AK8j15hKK42hKpY9cTleN1nTDeZ2sx1RH7dC0Z+E34ytVl7IRy
op9jAnsXBQDKTlVg67ziRRboQwqQ30/IpIwkGflr/RcJd5vNm8IfKBMKryR+Ogpu
03qHfzh0rETCIVIjK/pwJTNGGYhtJWEcKlSovChZYmgs4Hkor8MgoybC2DsPEMiX
hLL1WJuGnBaRTBXe8CJjRbE77WKe9sD5AZFQ8fIiy/vanWu+j8rn9/nbz6uvATPu
YwTJX7wiAj+jwN8cnEhkLD+ClvZZqsM+bQzUYbTxIfY7lId19s7G60k9jF6UtMR/
L4eUo4PcPuSYvzspvUs+ps6KLay3UOuIqUPyNvwJ4oiuyGKRS5F19OKvxQPTt/YI
u8R5jC9ewTnhoQaKVyCIM7iMU1DEUZLdYx0w5L4vsXC+uUM6DqNNywyX1GTqqwJP
z1QBjCDTMqae/PGOGLRjrY4aIBXLq2df4TMD2WClQEfI3zh1j+3nceQOeq0S75cs
3cL3A6RAQr59pzi+VeWDrTANsIPc9M6WSbSI03Oxp4LscxIw+x1W9qsJGgaHkVGB
5Njmkw/c0CK6jTtUGVyTsexPBiEuyMWUIHFUJkBmo08pyv18PW9fPPirnYdQs3pH
QzUsDTvWatlH2YvT2LoGIWnPcnjzXwr5JGKTz0ARkB8QdgXss767y7ueTetqh46N
NX+R75FhpxiQ6lJslMOluV16VOQR8FtCmXbEP3STk6TmzFnLUQxzzLUg8f+w21rS
TuM82NT7hGuY1sxCctGUSBl7uN2WvVa7zOa3AO7vk9qgndbNbHA+pK0YvLPyr3Nd
IETOSQer57oy9Fo0nwFwM2uRhNlkjezeiMNOf8okmPsD1lpvuRBP3x/DMFChAJoX
a9LgeWgDQXWJ/V20TzeuEtNZ3jdPXw5CNLBn5iPiH4pbE8QnbEfX5zuFOjOV72OY
PBRX6RB2hdQ5m2gDMgU1YdiL+DR6YPDVMIbwL6jWb08iUEx6rHKb8jBu347f0P4C
IesWumj8h1vwpQo3GOeXe6F2tFZ8ba9CcJXRSHdjMITyFk9d0XOYqIhl1wgSmlCV
GKVqKE2K+wppms1k64hS/tQNVWj85qpu1CaouaW/xlzo9GEoyFh+QKX6U/+VuqOZ
04RHseGjgPEbme9qmgz+gqf3Ze/snYXMtT9lqdGLOFstq5JfeNwfQLWb+K6iyV0P
CAjKDrBj9bBjqR5R+xxH1881OKih0nyujBjjsdIRKg7qSQ3WhOltSQJjL+hTdMUR
/cJTeMCpinBBODLyIz2yPui8FDuB3mbg5uugYPCLWfp7kjuTHFfFsxf4kLqFbolh
JD5aidsg6p/kfRN1snGuy+dBwldqNIWZAUQFYzsy4z9rb0Fz84WOQnsTa0mtMxwB
+dzjENZmvMj3I6owXbveK8xcrpviSZ64cXUjK25NFWSTm9EOyAw52Dn2Zx41AR7s
FTcbBuJpoeK9TedVOo829k/v4Lkd+85OTwH7RhZ1C13JmhB6T9aeapuqUJfhkXSV
m9VMbP60IbG4swk3IA+HTcpzOPx/JEVZnWIZn8BwbwBZYCsIR18QdyVzWp8zYdgD
Idc6SbS62HTHGo2+Ep2NF528uK5VMaSyNjNZyKZKoShpgQjPPy4/atojs+1rGexo
kTnCTf4sBrsnLTNO90ACo7UOOQHBcVPZyeWbLeHqfpedNpM3ruwIGk4j1tKpqQXL
n71d8CUq/Titno3m4FgZRaROkUFjh4NZvG40KcB9ssuITq1v+SCV3ErQQlMU2rwq
Nu0WMi7UEES1HtdMk6K+DksNJDZMhlpCiCIqlaQDRwVsrG2RpPAHyFuRomndnize
C8d8qo8AieekERCJGOtOtQiCyPl52fmo0X3tGhzxCdRqb6V7xSvKLkdMkyNyQMN0
2g8D0YFm8om76pcUY+I/1uJs1J44BQXc5bAo9WjlknUIg/gRLac012t8Xk91sKFz
AG95ptAjp7wmiZ7Y0cpvjZuYetmApr4VIp7VT0IIaTC3emuOONA/bUbpo7VuRSVQ
+FuQBajLius7Ql+ZbEIN9FU32yoWyNs7ajwiguSLTPuRYltjg6jcyi4N1xbHh2FN
K2mfDFV/Uza5gtVb1Yv6usHtY4tHYD0BfUZO35zVOvv4958Vq7YO1traNG4xDn1a
yU5WcR57yCE+CeJFNBbRemhWHTxm/BzyAZyHhCV9Y0SDrbSpX3Yc1501nMAi+Pmp
yuSExZPlvg+m2o0kZ2iLGlr+GI/3AeUKNv4UbEwO6CXNqLjuvS4ky/CfOKJIKO5L
N+R4duP44RgGJqkMZz8pZlHFx1MH802QAQ+LwQF7hdKPuk81h52Coik54IkTWggy
m51KZfAYxLPGsVb1sF2zO5BsPCW9o4+RC44zzt9C3ZGan1z0XVxQ1R0cxNxwpcCN
H1cZ/WY7SfjsPsUoa19ceekHYBC+1xo3xuSvD8oLQh7n/OZkSsHPCuINlWA+5wpM
x8Wanqr6myJOZMoCfSOHcYNsaG8JAJmSfJkNHss8W4zqgkYunq0uv7qjDFroWC7v
ownrYVNxykE86jksBYtppqpr3Nl04hRpEwMXR655ZcuNP/lwrNCpR/GyMIiUyzRp
hmZwN1t4jvr0eGourx9uNpKGJ9Fl1+wHa6oqgppQ2+x5Q5AtRmVm9RF2D2/762Vo
OyI4PPBUUUGLUJdrKAi2T54orh8K6yb/+dLduGN80zHO8gqxMZZsyU1lmrkcRSGG
X8rcqdkiC4qZytC+lJ12OdFYSD1n+hrHuXRP0zhzVxPFlX9Q9BA/cZkARdo1g4Js
+3s8GCZJkCChWb5xx2VarL8/JI5+GV9X+p4zVYEYeBNOqQ+PkLmFe91AQ32RfVH0
/UHccH2PwsQSNN8zAnBiX9h/gBE/Sp/Hygpm+v0qGzrXT3frrKuaQNBY6xKw4Zam
9f9EqIjK9/vEPIVCrQEbggy8YoYQl8jNms/E2Zl08w7TyrmbTUknHwRv40tg2wK9
CIFhp4hwz9H2qx7ojbB+N7D59l1HwHbP0PtbhkOCCtdG5L8OcaQAuI1hRgBIxq3+
Umxgerb5qf02uv9Znepgh88a4jqYQ7nIfPYPzV0URoCQ4JwYCuHxZjkkFOwXz9BE
zuwjl1SJ5ys/msI6LznLh733U3qY9tYbFexo/3W4P0e1zb3XfZMGR++TOpgwdV4w
C4M3IN9NXCcX5diudvIQU5x/gEpDEECPeJ7V19OhCWsl4EHws8o/rufRhYZLmqZl
3xB+0yiFXJTa7PrXzphDDuoPdlmtiF6YjgITwD1buNqPdA9l7e34HChBBAzWhnPu
V7ANSjRykr28UfUWhKaUUHUIWByyVajqHFPKyImpePDa3zokWA6XBAA4PATOdO/W
r9E3DnBPoDNvA05IrWHZ4hImdx8b6FsjhLGfaB2XW8zc2qPPb1rhoJfywl81MiZA
AdfwKtTtKF7tVNzybVDlbFEUmC972KiHTl6fHgROFXU9K/nE1hPSsBcw217tYZc0
rOsqYEkZtp1TR/cTQZ6Fn33WzYqz9nhuaG5SN6HbJavYGYbwonXitdRRuIIVRMM2
PbUnmPplcbpyswuZU93+Fkp5LDa5muhXLi7AEwy6OsVEfg7aAP+fmd770lBg6N1p
vbAdBXRYqgWPIUvRAYQ/NE2d3ZC4d0BET0Fd0s3b5B5kwLILJgK+rN05wIJ65urm
LH4pQhrZoLRXwszvRi5AlI3Ne5zDFvwmiIc+iw85WWsb/81hve1R7x41yM+v0C2E
6ZdDZWWy1ErrQOEcDEoBbwYVdHCnYjDchx5PCnd0xHd6PO16PTXukKRwB06ztrh1
xUxlVLuQK5/060NIKtwtontDq/hHNRJHI8YskaQaGjqHyJZSGseOn/jPD/Xditz5
a1vZn5nS1sTIcDL0qk2LKPvZxj7b9ILSXG8oD9l/a358exomJPDJz+mEiWjWGsg0
J96fsq3x7JRYiX5dduUv1UqjVks1M7GMcu1Sr+LwgV7ab7girz8pVnuv8iLGR1rk
ykx0iBJqF93IXOb9fVR75a1KJgWn1LdxxLol7Fh9uIg71LOevbkRWPYzLh/PFhHm
plUlWsnlkUvN+gXMtuc/SXd1SMnu0lj6NwN30s5izXvTye5A7VGJu/pGgniVWmMX
i3ciU+BkebH8L0nz6ZP4Ew7OWT/8j+pVcnzyt6Q8f4QnJhrOuKBEWxw0hfZSNm5J
BysUA1ci+3RG4E8cPx9LbujNXmcZ5baTD3SlBWy0NXUO7zFglwnsOWHPioEbqe6w
/7Wvbo2tR4bsSXBA3zINS/vg5e6E1Z5iVoZ+sEhaqc56A9gsG8StxE6K11n1KFzs
+1pzP1onUxasVu3cDT6sa16DR4VZZJ0x30GIm10B/3moKKNDjkglugAlK5YY4NER
ZMs9ST6lp2ey3HgtWZF0Bomdu8hDeaJR7/NpIJjU9d9pl/zLNrc0kzSsWlTXq//5
OJgEHGJtivSMWzF6YMEURxnkmrbAiQiQEKFVvE4pNaYBpMPAsRtJNY+7sDmzNCmI
lbmAUtX7fvbLKAFfUZjsyHuE9G3lBpPsU7TanyG+xF+UZvolqWHY7KqTmoanLyT4
cIzrd43ohaTnlCpjRMfeMB9YDbEDhP9bc91ozVL+biiSat8wv9OMv6VN2QUkvrRO
AXLyAIk1OogpgWUNIsPKKLzPy4gSraF6DhpFTsVsw/yoZshVDvocn5ci7EwYujyR
N790F44IRLlZeZk+dn36/KCtTJgCiHVKvFyvaX1iiq5OR/dKLy0nwUh/OGjPwLC6
b8Ent7f3NuRcWr/wmFUiUNnpuvRKQo6EwBUEBcN6XSjZYond5xurxcDQjqlBvdHB
UUkRFol0szJjciz2Tnog6z8LdIoAmVe7UFxalIN+w/9d+X9SeizFBL4gOyFN+H91
5bkmbzeZFXdsQMHFITPje0IcSBjmr78kVTKSyj3ykhf9F01+zmlP9XLHBtKt1qWm
/zHmKFwyfJqkFqdEzMKykAfKYZxxQ1cCdQ7K20dFT9mOJ29NtF98enjQl/Hbnoa5
+szlDkGI5M//MstHx7W1vzuabu+0cMiS0QbEMdqXFURnAjrOs5dzpcKzakcvToX7
jilF+j/6PGZ0gZX+K4dt7RaCofqHrn0QRCBKdEAuPd6bAG32cDd6rmm3NlT9SP1z
ZYvduYpIuZzEGND/tx7trwDa+ah6ad6Ze85hYbdrJhXipMA1Bn4P3GwtH2eytAWC
kaCQtf9RSBASptIoixFBuqoWTWPruvSaNn5Rji4ck5ZOqw9PQ/YNVPhvODi6MJwf
HC3Oy5M1xJnN6wZGU8LuByTE6frGf4mUJb8nC/CdXQsV90ZYLitspw+Md8vr0bMu
0c8sMnvORjPeFQqrHjbGTwOvvzkSrphaRgIGeNScr9lHA16iHJAaXbT3FEGDkhlH
oyazU2YFbC+AmE65vURWUfmxa/+wZ6D8PugX8ePNyhw+9O/fFxXjWNYyazQsi/TI
IKA90taDIYjK4wDyHL34Wl8QMN3uzZRJy2sb5jVo6FoO3yjy5Jkg45K1VnRsHph5
wZQ7Qe57Wx82SmQ77TNrSitWx2lxL6qpE+mkmwZtxCH1cjnO7RmpGAG68URWsFwU
vpTEqkaVPCcFX5qXrhwUy/yLRxPJxgDbeQ8sTNZos86zYLvVQMH2riryPqU721mT
Sorwl8SQkFBkmWRZaZBet3vTNfaFlSMYl/H5AZX8UCyfq0UrBnYNaIw0Z0KoMTTy
ukvzgX7fSjhCHJZhJYzt7rxajE/0jHklwSjWmIPh7JFWTRVv3XWedQYZbYeD8HZ0
cpTdj2U/cK9sAzc8cSVo5eivo4gNAw6LTdKWlo1BS8gUqvFqYxgtPfNHyh3Tj+l0
5IFWApIgZluU3LNYu6aoWOxDorIRzCIkwpsCgIAXi19DwOtqKzCnrJok+ZQyqe6G
sWm3JPdKuqGk1Wdj4gdhPXkTKg1QxsF1+DZIXqOwC1WV8lvg5robk4SLCzNjwF3R
HoVBsVbZnm+++7KM1JMRSJayv9Nqas7xg1E2hn/bjvDUHPbd+I28zWRO6mhMdwVO
mVxllnqc2uIniOX7i3Te4yz6mHtOckOUNeANv1cuPP2JE4NVpG64+5nrUqfZmMoQ
0OIQbbNEQuoEnnWrK9wHxA0iFcbo52pDVbWbZhioEduBkgdFAPhQvEi/Aaq4tbUD
UZn89WSGqRJ6Z2EUzncPavw0kslVtOPwnHgkFfpDwx+kmsMm3XGoLj8uX4kNZfrX
J6EphigJfFQ9DGdFlB/o0a2a200KKKRQ4DFgkFIeGsclzwHq3GQ9byeEMHPeJJLY
p2Kr90ou6zZwF38nFJAShBPaYDmmr7KA16tHRlwcyEfvO9Q9kfwYwEVe6DumC6OW
0j0ItQ6iK6hS37t99NP7QacJwIJjMSR7Ww9Yke8esczO0/LAKNeXASU3PSs1PQXc
NK0C/hUFgk5lkAu2gCMDVw3JS4JHP4LheTOdNJGdBpHUUH3lXAKQINB87E5UZOoz
uQFjUa9lXyJOPnveMy49GRoZXidl8DQab/G2Q6Zslx4I3KRMVUj8vZwjEUzxrBCC
PvdHXiGgG5YZaQ+tSxAWA7M6OXDQkZEM/JCTjxsAk1B02KSceDmr98XJtj4pOlOp
unt/WFj95PiPF+9OK8dUxgKBehnotWDKyrPvQaVKUSosvPZraHEqBCzeO3uHx/hD
5Ybu/8yI2wTc90AkOn2jWNPG/BWupGJCi+XoIgPxa/aVWpeMJK2fjdD9QhanH79H
Vw24phPd10sQjKy2Cf3bprQmRWHuhTAIgLi/wQMOvCCp/ZgqjdPfiCcVgK6vdHxK
7UQ9xHj17KU4p+ntRvndv/6eWsrh7CwfElrc7zRPA/Syk1/9aIPwkDDRrVG4gn+i
tRmfGm7lhGh3ciZmVCljFZKFKMv33DgmY85OxMKKa1maLfolS3qo8P3dqj8M5nrG
wDAE+FfbzD7IyDxpgpAw79AXLAGIgMBVvMey7Jq5r5M9WcboT3l46ueLOCdGlVmb
fKjiF1gmOHUw1QI3M9r2UpKQCaNeCb2nxAsu4fpTICjT1SewOwpoHkigqavQGshl
ZzunPthNMNnuSluOCDVCeRsf63FBa+H7vr7iA/H0ejd4asl6BfEZSEKoi08FAcyL
5mdgoHDpsnli3cB3wIMEGfTl/A5E/Exe3DLAiVv/FghY/G0fkBi+f5lchLPm1622
J4oMA/n2KUm26VcYalikKqymVMV+FLExIoviDIFXnxwZp9ssP8E2U4+ELeorA4Iv
M9UT3ChZigOzwZttAb7netA8ujM8cfKCwiIdbnZsPhmXg/woMerP1lPliLzUJ1tL
OWvp+pRJoVlz4h95JsuK6I0HSighSiNyDvhFwfOIrqBp9+m0r+vHhVxvMbYqTLC3
`pragma protect end_protected
