// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:38:01 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
cbyt/zhgCPOTt5OOhbJ4aa5KCZedaf+AVznXlwOMTBaoh77xELb+JGdjVL6Veeq8
fpyFaMf4Yj1tQHNOlHjPWml3IuwOiMMKufipo31lidff+PbhMDn//5jR6yNzo18p
B05x5oI/pRQUzUtB19RRFDuic+8eHENWYChnfS1w5UU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8240)
RJxGq92dm7EU9TI8XtaOqIDkhtKhRyRCHEGFBhNLRro9Ts7WKhoSehdDF86f+xA7
84uyl7JcU/4qUHKRDAdxT3/xUXcFyX+zMxnSQVXXcz+AQ0mFdVMH1AHKK51F5IAc
4fUuGXabkDmFPbgQcHeN9AjjdDzVIDuv3dmnEV+4N7IFyRiC0zHour/jVuufF4Ub
BI0x0FPCkpl+lR/br7Z7YecKr4HgUjMUegcqsFCXqUMf86SlCQyV2mLztsKNb+7R
kr4FxIOWXsfDGXHNFhnfkwsKj1oOmkRHjaLlN1ZgTzV4Kdvind1+1YX2WdaU+iiG
RkzCFS/oj/ZCiJAry7gDkSSs60nT5MAe81zzXemTzt2JN4MP52VG9NdneyNXi2wo
l4uQkAOSI2TjW14g20S93RAmm0wC7w0aEJBkASy9bFg1QcuHpfcNtM3aD7OtzDv3
2QJNjpmDfpPhdtkVh2nNYf/mXKm3FfX9CFcDwIEaibopiL1Qbhy1MHid9dUdXOW5
PT5Lol2Rk50AqjlfM7rnHiLuyN6e2fRa+MK3k7Y75mlHPkDnUOdCjzevobivVita
JjzZH/3gVRXbS5Iq1tKG/kErR9VZvv7t1SCCQQysNUjV67c/K2PASq/JXRrTzZTq
vD+8HyRUW5h3z9TKTljXgmCWC8pVLmSFQRzJ0rauYqTcY1HMKZOI/twrBonF+xBV
9jVnBEuSnkB+NmKytE0VQd5fVejJ6HJ++c5mEdafw1PtrTut+rEloq/H6iO0xR9q
TUQHdeGqZgzoeyV2fBMdK3E79T8wrusOTdyfWSbKJL6b8LomF2BmoROuC0rAwJuu
VFoMgnmyYwIw5IdcjnIObSXtjtvlJTIMbiqdCAO71hdi+ZEoVOTLu4nNq2oqd6wD
l6s+LWF9TotlsGoz0v8GCzwpbDgUbqRqo5mz0ZF4sjSdnEtvjYSemZY+vEC2Mkyj
aKm4GhKVDco92Sogmfqmg5E5F9615QgLuSoBWiCorj8NEo27BHa5tYvFAiddpIak
79BLYbC839nlosGfPNXf7L/g3+dzDDUyVvuc6uJe5VWK8vdg/vvw6FrJxyQg6HkL
fyq5P2ck8z4welgbZB771tVGehKTzmivA6jxddCLQyZc8YRydPiBhoAm8DHp+cfO
8S5yDZrvGjQ9AweaBeiHMlvZ3YPnLqq3Cm40yl+tFpiDcG1whGFJU2aaUukcQfKO
1hQVh1K02TXA6DvkPyBxVyMuGR878XxitMxBDjbkLhO5GjptfQgMueS9vW6KHK7O
iUIDy7vilhqa0tIgX0+uahiSI7c77t2+b6qqZ3/l3K0pkaAYe3RxTQrifuU4D9dk
IJNyUW+THuAh1GBdMcn0pThf1qq4mjilR2yIFLaYCoRaYU3o0o3qLK+PWTtxKvnL
tqT6PaZdrb10y3VA/Zva3vaoupGAjDKOk9XGpMXOTtvm94NuesZdMnphGuZHCVNe
u0CZN06hRW927lzZTDRjb264cOzzu+AfDN2xdVzeSGAVfUqBVV1HekC1SSn9fl5f
orgfMRKOhhu4s/VeCey3dv8HsXHC6aK2ucCUV0J32IhxvQ+SHJ6wAyNKnRyL2zhe
8M3Kh+FqmrMYign+giT315I466Hect+AuTTa/7ZVHDuZ6TmtcyhMs9dkzHdh+Fq5
zXNpYYKFBHFuHO42b5PiZBBGWaryYqtoN55JOQrYrOr3XbEg34C6V7UU3wcEwwZd
G09J98mdN+C5MBy/ufpmz5CbfPg0iQd8rB/0Me8HAzzPzdwfbGTZLmLWdLqTqwB0
jn+Hs7MGFG7XH7ob4oH4MZojYpSamsvXH64KxEufqgR2yHzS1HofEQai9esFGUsO
aIrT5YHmp+DtJe/FdBV3FB847SqmUtOU08/kvRGdQ/9NKm9KN2SEi+O5y1rrKHZg
VtDrT3gJpKyLFldaJx1qHXAVmN5C7yJIIvgLGtNcm6/uUouiXUbUfpZFY04bCNb7
GyTXuSkQDWjN2p3hfExtQ8nnPEPf4kgbUa5WNQkBpi9F++xNC0GlL51jlkVMNQbs
9HmgwkTNAptseBZhwFiEzxxm/+fETSKrK4yMxGH3nSN/FZGq5RbR0s3sOCO2ynvH
/ujCXjDBPSFtXOPr242Lz9fNMVJ8LFy5Ws9jp3a6qFtp5CMxD64D9N5gbSJrSJ6l
0LFnCX/NzErEwzxWBtm8v87CPtzMEif98gj1UGGhDez+1tc3GEbEey0W1zWKEZZc
2ZUwco9zRQfCt0QrFVxOySt1aREXetR5HcyTqZs2XxuXNjSiruU43EqGrnNQHoN8
QEHa3vGKMO5x6H8HlurXUiiOIxAwrQa2ckMDx0qpb5n74v6ozlA7EbFRBxWE0KGV
88MOWPXjSKVJAmBv2fNhX7C++DivPJjj8Es/6OFO9jZWhJHKTS0ANhl3f9Vs13uC
YSm+a6JH7PIayUlYjYAAuVT7bNn5sQSC7FHdd+hVVRfN337Qt4TAmNglX+193/h/
lp3K0Ou5bjoAYCKhypKlqUHZ9mtXQzPqqHDDD4vJc5bEV+9/17MM4rg2kRBp+pDO
NKFkdvuKZL4dhpsKScRL2sWBBzrwB4OudjOHtDx246FJwiFlYg69wKawZLPOs0dx
52I+BqUXXm+CZbgWLpB/j439saoeYaFs08ITH3ee1MUTH4tZNhBcesgmnEImhQiF
8vmpKXtmJFH1qZF5J5IqXmFDXxY9wxPzAwvn0xeGbKHh39tyLrklKFzbCI8vF19Y
TtZNmMyGT/aYI6Bv961jU7nv6s9Womz/Dhh2fVp9/nV/uhRU1iS/12mlhKFMEOkX
Bc/2/p9DzB/CXhGbnfC+th4O9yds51a90VEfe1dnkqe6JhuLgMB1mI+6dIJ6Of8J
ksg9PyfbptkB1MmN3MK7QOluJMXOIE/KB2Niu/CsNI7M/ItTIsjIw10brgu4KDxR
NGnQTPX2zDwgbM9U2bTemhR+1JNv4TYTt2Psh4RNTS7hdQIAX99/h6vH5AxFLL3a
UdMKHJwMUYSe2GkdWFP1pwrHxI53JDFFGgduIIIrJ3CNsmpkpKURLrqr2g3FpjV0
flam0xlIixY9lVBz6xSfNrMVZfEA7HHsBozCcySEAq4l0FxQG0D7JAfKWvHH9gTm
dUc6bHtq1YDp8JB2pRxPlGLuGeDIt/wCIseUyuqyLXQmRg2ZUo4bU5OVHVE48HhQ
KJP5+YOzlq96mptd9PC9bsdkftDzihAT31kkNq19rAJl7hw1GTmi2zszw0K23Slq
N710gwwpo0k92N4q4sgvWSCFLdpYTRMsYq60Ym5u4VrGFEQ3hvjnWtgGKcw7v5/s
xIJpLoCYhFELjDuDbh3VI1H8HOxBE843+joxiZjOF+rGuK5E5mK3g4EWFFu8OVwu
2UXMW6FlBldcu3xWLXlAiPUral0k7n2oJ7iihTlalqCI7tJic82tRADlXW9RypDh
jJwE+a+BB7xYJOypsHBzISr2y0a7bdhWloEBqtLmpP8qdmUwThkESkL7Ph2ko/Ji
tlvAzCmkFLbcIO2yTh2iv8gCYl6YzpQkA1/UMHP+AW2p+t0UYAIA9PbGwNNV0Z74
2WmE63vqJIC04VDn+8xxrgIhOR3HktpD4stuZ4dkRCrEJyE6D0z6CTvzh/fAFCXt
D1iqIkEg+X+e6eJ3hXP0SEBXQD+5k0LB4GNtkAWkRAPYc7lTtpBDJO6BEhX8led5
ZZqpt4M6jupgUkm25/O+Wrg1bp2VJ0+QZVLHBPK7o57tDNvB08C5rpDHO9Tpkuqv
PQhsltSe0FPDNNfGoQtSCPyoV64mw2g+zziTlNhTKIi+bZA++vhuGBbe/zPRmrFl
PZETe7ZO6ynzBpguHrCIfzOOug9J2rxlXDmm6uOmOlAY7T/2bQGBTcxmcavMIU9k
QakE/p/+2fhwBnBv+weY+0+8mF/wZ12lBSZLuz7dACspx0IbjhCn4MtDYtgtJfvS
N4YINdGnCn6A25bi/YjI4sMprAYi/0VUx7q9TrfvKGJtAtrxyMipmEymvUzZ2Sgt
fhZv1HaxmG1YNFEok/RM0sGA06IEJN/WfrDa7XjY/x/bgn9wFJsYMPCERKMVadVb
LNtIiOaiiKhjnEkDwBhMoiqehRnnhSmbPjX6kx/Nf1yl9hMy27ALYCLTcY/xxSW5
+jh1Yil5ucMXJ+ILJL9YqVH6AegQIZDxFsALJF6akLUg2/h7dPMA9cJpFMKobE67
tyWYEH3b17yxPmSxTmt+ng4ib9sg1YBo5bVX+95/00YqI0WRkauXxLwC2jd+HdkH
44khSeyQZa+IGbvJ2eQdvaH29Lr+j6JoxndU9OJAra9HIIOpNl/lAO/3mHAHoSyi
jKwXlKZhlfuagDoer7dzEnciBblqQdAI0vVmQuHUi4lV8oT74n0STTYftw896WsO
nVkRDnw2vQPd6N6xWsekJggdLoN7LCSu2ZmfCgMlZlw4B4V2KSEi6bEpXl5KGwQ/
hGOWHFPUiCOi/6Nut8Zd6ebfV4O2+t3BlwO7PvKyWCHsxnaLLUfcw2xGpXZR/e34
0Ytt49PCuZBviBrLK3gc5V828cTpxznvKhE6cesqyGA5ekyxK7WZN0vihWlgNIzd
1YoGB8j60ek8hjpKGMAF1/ZKNC8dlDOP4zM03k/X6eu3zYO6ZNsgFvudaHoOBvgB
B30DrMPEyB0ikJUkn4TSVG33Fd/63pnjNIRDbdXbz1F7iAlnRQnsx++AcnLJc5jQ
42eqIRVcEDFX5PxAGoMM8G2cOWDeBGt2L1TiDE4UidtmsRBo+AtvcegtVIcEu9d/
yO2PjDtNtt1/B14Z5P6gc2FeDbh+X77iEVmtmajQFsTL32JQ8nNORrZMxoZs2oLh
fn4mhjNrhIxJ0vk5gaADG0tK+pmv6A+XWBMBLybZBgjI+rEEZfBVCeU47hAUQgW7
U5823ZfvBiySY75ubLohBfPKffVa4IuWRrsXQg3C2RwpvMNPhjXRdGL7lPNsvx2G
2iV8LYg30W6fk9Aii63eAaUebHyVqgr8b6HOYn+yg8DCOroF2YXdmOOoMVDRxK6L
GnJeRHdfeEzrRcJzWbcoUW0LGNQeV3dYPfi23fJ7IWNiT1UDl+ha8OEdYcmjykBG
Pc8B89HrVbQxO3y5QEXfqivxvTIhHZ6xKFyTiKKfLdTw3XgX3dewpCgHvrIA2yNd
9leR/ug1LLJUt7a4ZlTCV4T4whgu9o92NlBilsVenH/3pvaNZ5XpHH/8WzJHlJnT
uuFO21Mee/XpZKbkfeliPB0E32YznehtDVMDQFuC7XK7coCBXMyJUYoc5//dZTbj
rTUuKsBClkN9SDMmH0Bs4WaGCnooQG4Spx9EH9p4wEoZ4BRgbyhCdNO+GTES49Ee
TyXrd2UvUi2qXZR26RNrs5NxU5X61pjfY7YhjZZMajqKu5CGi/7Jj+83q0q/hS66
2j9el1qBmtWxBfwZ4lIROPQzC90k7+Jgg+ySmQDtr4U2rEeEeOXqFCrGl6NvWGIC
LFOqB5csVQtqOpcL7vEOrAyAW04BiGjOnS5aa8drMrbI/JKGIFmJ8DS1EQYmXZVX
CmX/twu3Tfh2+FPWWdmYh6vmrd+iTVMBseEANzGL9orETp6Ztiz+un5PcMADsEWN
K+GOKhdOW8Y1qOyYyBypHlrcUPW1HZxr8ZsfJ+JefbI99HeH87UWH0HZ7N4GcVh1
ZmEi5QQQBkY4KUo0vrIbgB9TmO3hzIRZX19xWjcoYsJdioVFDEHv2MoGsvwTaM5H
uqKvUjHZvXBoOwxlv2uVj3/FY4bmDrBujrceEbXbU8TvUaEAkTTQ4oDwTEKeSlUw
EHVSd/1M7uiWbw3y/vM6RpKJTfHZPGyabj9vpJ0B2gcXcGhWrQQ9pSiQn6HS3FUV
FyQzSCt6NQl2C3WcFf65EvuAaxfBy5ZNiKBGFcO20Hd+64efiGdUpM2RYC/iSjQv
UrJOZaod0Y0iWnWYPInUqqQczfLhECKEQSKLj56MnXWmApQ1mWiJrDXVQygj3pDt
hOz37lNZYCZDFFN4EoTFf80+kpmyxrIbLfnY4+srRpuF8ehR0JKjYgLzHUxwc6c0
rrtQRSi8zxoE7L9OHQYgBqPj95lQTJibIYzteRXBEqlZ9TTZ2BE1cjuji0IzPIxj
GB4T55DFqbjdNzHj+FRAUWUuJRhjAioBO3Wkd7ZThbPpcfi5LqTMUnJnPcgHq0xI
lkyPGOpgbym9EEkL86HLg/5ek641r2b0UPn7e4TJVO4BqsBSohMi3zT8k8bE6m/c
AU8F01zDqnSHKfNGDs31fVlH2+rXslODE1UY5nGJT/jDMrWpoB7Ui9Ug8cskAoiN
n9GTKmWeBbDZQAOS6zx7YPdM4/XYYk5uX/4nFOYAA5Jfhh8u6oC+l+uxsKEC7y/3
z3UGXh0wa42XwcQv63hgG8EYE5mYTMtGQDZ2MPPw9bkTDdiKt0yhT/XhNX1D1SRx
doQsRiui9VA55MZ9AS4YJAFf/x941ixkU6NEbvS6+DMKaQ2C7R6cRwl+CZ4ic6+n
6UHDgfaZS+gDvJqAgdb8iXsH1JibPxsFp1UZ1DVlSjMBUIC3LP47CrfrZnIgO6YT
n1jrHfYy2fwDN2O6GhukrD2tji5DjCg6ocoOqfOWK1DCrSBmMEdJpHf08T0T9xee
HCIJbNNEgs9SeG7MlpYBEZemn08sCcFRCRcVSdFz7MSUF/y03K57VxmAOoBRJ9kz
uVrSK6odokPJxRwZBvcmZfgnuJhibpB++e9rrGzixWLM++Aj/b2/h/oKhXtZlrLQ
jKS6ITdlglp42ZQB6HtXXKgp6ddAGgvbyjgEhMs68VIvuEgxCziGlvk+FJZvjKwT
Hy49g/am8JYhM9+G/SdT5B6nXZJX3r1uw8GiJBJ2X6qDdv55TtBs/8ZtTOVPWXCs
A3a1sBJ7wGDlX9MyBupZv5/Qg9UWrZtUG5OrUDJ+utneeR9Y7oSkqo9mr2CXmFVt
DgVHUZyDJDUeQxOOyGxf0n0jWlUxEtMPlPsud7BCyQ1/Y613d93SgT7pGwheDLtM
jxuQS2Nkv9AHfguzmYtnVmuJVZLKpOk89XwlGYcHKt8nZVXMax6O9U2wSwqR1CPI
X6xPH2xCwYLZQEi+7ZHXmSStPqKsUVAh9WfZDVXP9rCIq2g9CnzzCYZo/kmf4W8k
vm50v7F7MvS0McyCcxYpqduAdf4QUjqIEfsAgl6LmlIbVpGh93GPfu+QQEouSZD/
/GyM5Pn5l1gDyNgTZT/KFkq8jarzI0dDFGHKUYLL4br3FbNR3UFYgsZp0pEw5McD
ESvG77N4lREkrPGgz5auYGbdUdGA5vcoJRbhHawtHLbPPaZRJtpIx6nM0PGAslBK
9s47OBTtfkteDrDlN8MpMBto3q/j2bcpl85m2OnTQU97wQKskBr9qfCvmAC3aRAi
BCiMYPhMah5tPKaOnC3ean78g2RAyq+oz9gWguRtgXv0Nfj/a4vc9okr2Hb6T189
grPv51x+gPzhj/mR9IEWQr9LB4gC73SAv89XCl6wqDU1aAd5gFYZ20WSa7rkwp1r
Oh1aaRU1aywfHlMw++cT02bZwtvoqRxEx6QE4LU/iOHql0ZExZvSbbspn+D3nXkr
H4Ajco6/SiwylIg121s3Lb/m8v0i3U8vl0Qs1Eb5pIIMUTglsR4yAQdKBgvL9eef
7qzJ34+gJJ3tdPyt5Xp+pcMlLoqaEY6xzcNGQiJZdhl/PC6ycXGeP8BGYBO6uxu3
s0w+xtoXm3HViOmV8o2gmeDVaOZkvIU95hr842161R4ddJH9OW0SPJ9AqtJfNwdj
yTEGCv7E8DQm5JPqwKm7tTTlfzJKPvKuKo/XpPJ3Osu8iuVJeze2SR+jJ6aC7uPz
JfRMy6yBrX8TDcxGICSeZIxaFR3vVFPzGfBQv1V5QPpMoqTXCyXpAhHTFVGmg1W9
YXAHkpVhp9QmYp9qnt8yUw42I7xDdECq7eXm251agvv5pUZUFY+Mql9L6VOkGS7E
5R+dbUrzLGTIcw5kEU9dhy5gA1Iesp8Sh+GOtkG3K026cGl1GVDYdVMhKdY3f/FW
eAavtd7hlIf3LVFTda2N700RvmNNpdIDBvIU22UjVFUHdQkFbqhHpJOPt9sJUIXF
FksuT5L7iR9OdTErkTbFiwaJffM9GtsJNSFDMSLCrFuaZlGB82vYO1cwI2rxQV2h
hs1Lt+J1blhSWl9lSsBzD+xYk3Dhdw7IHmroFBQ9TIDM1nMT8lT209iEC8Juk5bA
BQeRV1A1c8LPAsue4/IGnn4mQ1sNU+lftusFpGJYAWdiLhuYOeyKEmhDGZ+N5bvO
7ips7anzveumalvaV4qqdPYjwq656uBMuEzwjB/xJxjY2emnngDv4XF0n5cKbkka
kf1yquCLnCDhjne7jK2bcpaAqC/rkxiR47zBFLzdLFkKRdvbG7ZMXgnGn61Yyr8V
+D/xdxukYniIwsZzOoazUo+dc7e+T4YlP1y/fqixx9idisLQI5U5iHYAeOo+VArO
jGWmpHSKfGosLCJgOWa1YEJ2GFs0JVupLl6Qd09ac/vxFM6Ng1pAnmuR2UiuzVS1
H5qXIm2chwzu+Lt6DoM0Mh61ePmCc4QTFvXjM1bqJxfJdpNi10O5BdyP5vQ7N1gi
O2VYQJi2SYVO6AqajR+l5XvmOJDl6GYYrBqS98CZ9tdm5ABOz0/5vathmY4V+h2Y
2egIOGHj7ua4/2LwZ1UcAjuFAOoHUhwzv4N3QJGka5BdVu29IDbDFlLXYztZh4Ei
zffvP1FmsRUM++w3ZDS3X1hZhG3ym7Gpp1BMaW6GtHfU7LDLKZwB3hJ7S/JYnCzj
yICt3FZKwQDUOcSR2jn8M9iWx5FFczIwnF9sIksUkZzQtr47zge0+L68uh8/qPlU
d8HZgG0LqUpgqisDud+QCj+FRGgdBfpEc+bUHPbg72EAfmtVq29KMS/YpNOIO+q3
7Uso0cQ7VlfvF3vMw5zAd6HK7/c/3oYLGJGW31B2qbn3NmEU3RzBjHFwckC54shK
pxCQHZJJQL+DlDk/0muwh+HbIIqC/RGwsb1kSiFzQMSvh0f02GUHC0Nop93ipIYV
h3nG3CPUUTcXUMdchTs1BcDBwSzyZiZ6A9PLQRFHt9vDHQjqv2WlKYOd1aLDf65C
Rg3gmKigkcmMIo/dZFhbLOspTJU0E96wpzx8sTy1d4WIhT9P1IqFzOmc1ZlNZTki
/6Mm8UwfDx52vWY3QOHeRUaiOCPnMmUlers4yPnPKekMeVW52xmhhKIfEgaUILDJ
l7rbHyNRbHTiO6+RD+osrGx/u038dn/Mr7z2vDYMQZyw3wjVAPezV1I/Ro3/9FeL
CiPv6Q5aGx2oP8hWs+bo1DMSCjCsFn+FTOYcVE30HwH50FmlM1cqf/yh/dhjHdLx
sjDZQrt5Bjps7AFQXcaH49im5fGaO2p14FjZjE7gAGKCHxIpvT3kedRTPKgUvoMw
EgMrulakBHG1/0y+BummnVspdS09t2r8uRrBHg0c8bPr6s6pWvgF2si+Gm+x7szN
N6yGgz6mBDS8cRPuSrDViT81iIc4lNRPuM6jUdHO2EzW0OxFns34evlrgx35j4Bn
fcGgigXZjbabCsVaYdzn9kyq4sDLVbFNVsA7yKvb8Q+hMJU20mIRbB3DsuT4nRP9
g4q1I6yg14wVTXCyDNvkSXOczsA6s/y9huqfhBL+okSZS6232qR2V15hEyyOF3sd
qfyNynCoSLKnqamWAw2g0pzkU4WDAg7WNMUEH+1kQBCla4fxse6C+/chQBCXNn3Q
8qdYUSRycGDCHjFskQGGXaY8j3GRdrDnCyHgO3Va7RMww9LYhlvrqpt4D3dIq7jZ
/IT9HI9ygTQEx6hiMFUqcS25GZ5qdEP/lVXyz29wE7KcDx56IrkWs0dvoLDIRQ+r
QjsRJra75eMLjByClGhXmdv1ZP45I5DrisisuFTUulrEtfRK9iTIuvSP+n5pO57a
LdCzLaHHqlER06vkw6MHTEH4OtTOj1XwNS+QvsmfoxUlyVk8FHp01OahAZ/izUvJ
p4HEcyBNmRrT71jIPGEJX3mf9hLw/fM887+S8sIGQ2qGqmt5bFCdtMk7FXLEsYpI
wulBTQHR3Aqxu0HwKRrg3iDDZPYgb+uxkyeOVWYiIlXdrQ6H0/UbT9FypGW2w5Mk
Ki2uhrtiUUPM2y4DayfI/pobgtEbeVwUCaNWsH7Si3/kBD9LciuaHIOmdhvutxX2
dsq3e2mpg3mDR9MP/ySnvsnLBx4D0pJomNDABqdkANbAEw3Zv7mgxwcvf0VDvId1
P4gaCfdMvUHJWYFQhJDbsaamQGKc79Iarg7P0+Yl5fdQwQ9RuI55sOGW77yINyOV
hJXW6f9CrzuVDEPptOrIeG3UHzBgsPvS3z1sKmiQfXA8WF5r5W5B6N3Bvtiddie3
V9dqeaFvbha0JridVsXkDx6BJShZMkAeaBHUIWIindI5RwtNcWg2ujNbfSJjL6ig
Gyg8XE4YJG2gdiF+g0WezP92KANXov7YqALtgg9S64Gc1AX9MAgVB4uzT2CbBVEP
q0T4WryO9eADAu4VsWcmkO5otNbC8gD+P0ikBJ8HCzZ/UUrDoeMctCn0YQUhQcLw
LfXe9a0k0/7WaAaXUhIzy5l9bMTWinUuStQAJLKTD4JEwkVdlrW3gND0hve3uP3Z
5emTk778EdSR65Xou2F7N0nDWjmvc0MQg9tlxJYpQ/J4BRYS4iPnd4S2rpQWh5AA
coEA67KFl50ttyuMi40JSVmla4VdVWWNEO0xe66+xpLkc+VFxmCbcQzGLkYlOD/m
SZUMzOgbqfoTKvppDMHnTnGKsDf7AvIuR9zVvpJdr8CwPF8RhTl5Eu2EDr7GIRaQ
x3ANnWTcJdpqWewYSuRVMEkmf02vlDNrjpzNjdKY4Rg+NxC3W5W7DDZfEss4qqbg
lKejvDB68CARzJvZssrZFdWb/vDqFKzje3/ejk7iJfg=
`pragma protect end_protected
