// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:43 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
nbwe0RNo8NKHV8+dnD0R9EcPPRpddjz6oTHLHL1kUo3A27hNbshcwmSYk1ufplMF
4n8NbRL3Us5XyAi3Xa+UqjDP92leRkzg3B6oXzMcO753PIXCgBroj7LX6Hotg4JX
3DBc/1MpacMb3vVLKVkrHp+YWEJiYqjLyHgZ7HAWvd8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5936)
H7AocDRe63ltExEWrqKX7npntn9mnQoAILgyc3rRq2B2AkV6aLycqsE7IflcEmCL
q8dORMsbJuCdUL5z2IlhbgCbQ8FlNbaRXugxmXNQtVVi4ntgf/ClaANgB9ShRxin
qxk3KHnL2wMBTPcyqV/rEkU9i+0Fn5B5NgzC+0fVDH3nSpF2a+yTJuPY2KfPDyPa
HJoATKkOnfYKXyG5hrsuwb/75ls/BSmdUGMcu0XZ3CkHzepDHgDjj/CalJSmlAo0
TmXQS5M+PujYRvk5ZK8b0X5VkrQ+SnExyEocKpAgYULuxb1NJneiuuuvhutS1vBF
PTV67805yMR6gfT3R2Aa7LtmMMfVH5i1E1hw/tNgBFUdYtrnDa21vf9uaNhSWkkB
ibxOFWNv5LiceklNo4HybHaP/buaO1ShXtHpN9kDzJ94WJBsT6UyC0yuK6XH3U5p
3NVmOHiOZtkw0r3nMNdgudhGWv+EBhuJvgi3LBX1vfacbZ5ezozJ9fmWi6Rrs5n3
CD4kw4v5+901cLYKzk+Q+YgFUO0bO8hI0pMqf8dKzFljUQg7NYPKBXTkb1PhnSlr
cWeRvfLjZKxjlVwnytWSIBxVOVEeIbOhyxqZiwRz9Vr7Ws15nDbBVWlnXvEQM/fd
k6wV52sID/K98yICQka615FzfuWmkyjQj5eA30sKEIVQHfEGCLUcRdPv/OPeFZMM
1q6l4yHxXrj9dsgZPGf0ERJKPMituKwkTMJK4MRka3M2pmyl3e0kyDHoeWmmTYhw
capVd8CK8mHvBWjeS0WuK6p7CVpx6dVSOa0DYq7UtUj4hlmQAtwucbrfjJkXMx3j
Jhb311dBg6t4v3p+s30z6V0xh8pGeb25FJ9mhERYKrTnCKuaUM3upou6AdnEqE6Y
ZY+89wBmFY7FIbUJnVuDJR+Od4CGUIy9NNZmhPl7gkqMK9dvz+pq8p/iU3qD2DFe
BOG2XPrqV5bI+iL3Iit+t7p2McMrYAztxmEecKz/TgF2jcxUJ/PhE/R+I5w/yBDS
QwCrW5Qxf++59KKMLgbBZYzBP9+1ZelO0/7iuKKrhgpv2yM10exHH6M0Kcz1/J1C
CJC5hA3HEGNw2L4rgcMLwlC6dmIYdDoSR9I/yKqzMTTeoNHRAPS0fZcIqiKDwnZf
gdjanKkY8/+SsEbxvvVqHwiKw2nm5M/JyCmZxNVXkSyPqJcljcCLSAFavhm2aK0r
PqNn7z/Pw4bJDpm1XfZc3ygMPydObYyc1D/GY33f9dvMJGgq9cC8/mOEZNJzu8ZS
CtwiMmbnVqXPc+xxwbzy3N/SihZ1Je9GZcyUkWydTID0xgB+E6g6ASGjoGpji0rd
ncVIwjF2QGjnjfuKXCzAebGMttV2AvvZaRF2bK8panC69u6ARW0hcf7b6Zl8akvl
mHHU+YhqqTo72KvN877/xTqwH1jRnojPdK0/T0rpt8uL2JRz7NNl9BMMZ2YNtju3
1Jo8NNNAbtAuDDt8XSzyP+Y04z4uk+uuLQFDuI87ctZI6SA3edNVayPUXbJQkHIU
xcxf5TZtPIHrt7prdEToNc+6SxUxH++7FxSrU8iF5Uvi/mutK1fJH25V1SOR7JIn
5HMRYDss7NwVTwSWS3b9tm8RtvTAjDnEkx4Ilcewb3O7/kqwEwHoy9xI+uKPYQkH
qs3wh8U3XDNj4a78iydeTmPTmcpGjCpMYXup0dJUBCZkJC8efRvQPqSaiglqCmLH
WrTWlBN1CL1POBMa4IMSGXp8Io0JDx+K1iAPOMjt6rsSMOUmr8sph/UgQ2iiNg3P
Wt2UXv3jYuAVengmX4CYWnFtusvjIwuLGtTsm8dkbJ0PlczS5MPA6JeD7omsJf4c
6WpOM3ZSH0Ef2RVj5svekmgHEwB7C4nfVkCGd3L/Bz4MOO3v+34QFGBmz/O7OKjf
foWU9lGlxNW3z0bcONlAEGkraDTkE/ejp+40RGomlyTM6a4cepBJSmI8i2f05td1
crk0FB7jF7kl3EWNG8JEI9g63ZEc9eKz+T6LaQ2ffDA+5FA9oeRAUs3jtGvn8fcb
vJYMjY8DdwDzSR576C1aoMVd+r/VqeP3BHsJwG6r+CbCBqX6AIW1TVKw94/NSsHX
JcK2jWsnkVZqBOBtroQD9iWzwcgyEMqnPQqsrUFpP9mhm1sUUmcMogwnbqt4Ujyr
K8qtgUOmVfWon9nSjviyHlnGN4pyPGbEZyiKTqtTPXTCBMXT9uD5oFLj7rgloW7v
8r6FtqkbtjrbtrEll6Oq3rLdGcnQMrQRLoRn1dZ5g5DVQJxk430uGfupCfIXLOBT
2naVcJzEM1NfUzz/tB+HYLsv/E2DTcunbPqn2iFX2iyKQlwARXXp/8C1qbJhlbI7
iJFTzz6cDdaWN/fanPNEQJzsFWeDl8k4DMOq0xB9lx9mfRhVaPnnbyrMFWyu6PZg
y21szKEoA9+piyKdSQPASu5/SrURuGG/CS2drSb1/XBzlnEnf9FgZJv8wdxE2EK2
lB27XSpFhb2HTTMmHhptYfuPxmKyZSYe10addOTirCz5PaQHxIz18uSCiOtTKrac
Xanz0cSvRqslUCu2QONkTsE4RFV748mV5PahDOHPYy9rFI0UfS1Q4qrhGMT5aM9b
M5rEiuM1zvdXaAzuhs7zHcRE5N042JUC7t8PFozVHLoIC2iP8oxZRP7v7rJm9PHA
2DDRzfCRLtJgtwLcqvOfhqLs8nqbtD1OiurcwdmbtECkwjUx1NFTSgbn7sB+HlpS
dVUUKm7RN9cmKJ6scGv8DKl3buuGfTgXQ4BkiZmFx8W0ckzt8w+3LKmEII6yHoSW
y7mgdaZ/cYeFpm0noNoCb8CCOg6Na9CKk+GNbby5/3Q6Hxu1YhZbhndBrk1kBQ7z
ktz6+Ok2P3Y0XxIQUpZVvWNk6/W5xy4sS9/VVOX8sIwmxdaK6zICajevoRsmeDMp
ftRSiW55lkR9w2CQkWDytM2Vgla8W0FmyDc28x/gqeJnFb9TO2qk0vNGKkdJJVpn
JjHsam5YxR52ATqK+yoiJT9Wr8UGm0FzFklprf41GSDCf9oCIv4R4Wo94SkZQ1fl
S+jyPrvCEkgDIOE7PGGwYCnycbbSp7JMcOf04CUhCA/JUvvm1Jl9BK6qmVu0cqq7
OGmyrUdHR0Pz3GyMhGXE91IJImxBF1lHlWGp3uyLvChd2gcvq5X56bhcUZ6+BkE8
s25ZQdUOWMgtQ+6nmH5xzAn5naVAH6B/c0NiHaIdt30qGmkf5hoVFxjpEXmQFhnA
xCwe9LtcB1chFoSyzz2AuaNv+2kupBtMlfdmWpm0YSyxE61YELgPTGXfIzZ6HErB
U7b77Y1BkRIn2N9MU++H16bVi7KS38v+vm8LkxtmabW2gfyVRhqLhXVFcwpYgNWM
5zP3hciQXEf5MRJ2gR3y4cCiYwIUaJiBCUSqqL4wQBoKiBir+/4tzQ9gWn4v32Du
R5Ez+3x4aHbOOXJ+j2TjQofm6LUZU7igWw3CjxbhNkpg8AAQ4IvY3OKXr8s4q186
5YSzP3wIzg3YEmI57AK/Tztx62MG06SGc6FJ2fMTapGcUyYvtzQGHq2qPCZ4Fa++
ushcJSHf0WjSevJPUfFEPw6g3NTHWXwypa7xmSqetgTyvN1I+UyvRLmtRg6R2SUi
glN9a2baZXNA7T9eqZmTvCCFXkk0OCDM+sqcR3qTDf2LRFiRRI00+u9jwd71dgH8
/6SQ6SieaIFErSrgzDxdx1TJ6HT0b2ox3ZFnndjsg9odYONs0pkpcaB23aVSUT5Z
ovJ6F0yb+0A42lUfL4U9UTH+nii2vjUgYn2ALtVGEMUlx0LwtFgxxT3YIRooVvKU
pllbtxI0bTVDH5n69GsjufPy2SHgt8ajdUm2D1YQUcLXSaPCY6giPtWWsRAZmlq9
g15XjntFLud0/QxR988JmzTf5rq9Em/wUAsn+wM+Agx/90tlLW9f2F0CQWgwso28
X04pS8XofludjlRjlMHhws9L5Odqlg9s0GdiHbhZ11u5upAMWXZsqnCjPWBySNOe
FdEkCmS78T5ekhM2uNve3pWdQ6K81aIEEzKDBjY6P5MN1j1iJqI4exjLjoD3xuhL
OKEMZWA1iltLP3qrNWGaLr9kKB690gg1ofSNs+XOsY6ohIsLtuYzUfKyTxtNAopT
tJnPRIGK3IgImfAA+zwbOJz2LK5FAVkOaBgQXBtKqTR8VLtZ0Guxwx1QgvE420Mm
hxe+oEJ38C543ZL0rAHZBev1LU9OvMwIHZJLx5MbH2IFyCHkJppcN/d+CJBQNGsW
JsfdUZKajgXamyeLGZg4eg3t79B3EUECBXwyy6JKmiSRDrnJkmnDqb3zKjy9M8Ms
s68u2UJYtnFERdF42RRiNHPfmWUvaUktYhaUpegeD3A/+TtA/ue9AqkgcVdSU57K
4rtgGcOE9Zs/VBzus4xm851DCShwWdmCTsxjWhex6bNlE+KDhMIKBbZCMPwK9sIu
Sknp9JI/xtkHk14QolOnZr9Gywjho6m8oZayNfoRJTeuGLkso+21PZ6Mn2bY45PQ
X5TzI5oc9pfHZjmwKLBwy5mifR/kQPHCtDy++P6qkZZLlXeyxsC/uPqrk54X6H60
yXcIXfeHGoYEkA0a+EtEvGZyUQF2Zw0m3dfFOwqjUKByk6VOptNjby+q/pnWNe11
61TKkf2EviGyqgnxaUN5emstpZHeHC32GHaGpW2Xk9c1ElHkkxrD3Tw0knaT8/iU
HD+eH6iALVkUIQ6RP0VIyIOjBBd5yYz0KB1O1UPBVckhQmONlYzLZbzib0RRa1JV
nn5X96GjJkXhhB5zh5ymk3nSVhD7QHDe4fMO6QPliY+gBufCVa2NLmKXgW3zJyUo
PYOJJ6FAEiL6NOiXiehMIa7U8hQhsP3PQMBKqK80Okzy2uU2ABscIOIm2Yw5NaW7
sgujS7crY3ulCvuZZ4QI9ntjxIrDDfPTjkMSat69WssruJqnukubAwKnMlfr8ZWL
inK4VtrZ8KVBEpixBZ6gtZEdlSJ9pak1OuTRdVi/xiPCMxBE1BJusvbPlc8kLbBv
KMDhdqSkw/67AgrtDQTc59yMeE5DCRNpocwKx4drr9TyNzPLQ+HPVFRGDZoNLm9J
Sutnjz/BglZnLSK9FTOJa/jzFd6OLY+wNfDHHyTyVVPrW1d7mlZGH1SQaTMwSlB6
5LHCwz5Q57gfg/yWRAF1wXw/yzIGl0/S3S2ycX9gbiMNzn4tKcU5jJE5dZguM9Ep
69Mvvlm0tTtBeAOuqgQ7WxjgCJMSaSRkRsuKSKwdubjr/f2sInnOEFgDOeXaRckX
vItp9ZY8858puoqN5boU9fA9sGSO1CiBkf6Xw/ABGMK63ctUb+SfjIIzF9WiN/Fq
Q8azhnf8sL5IRUw8UiVbm6g9WcKtz8VYQsRc6fImS5w+SJXtKtOvouuf276SnS8C
R9xkefD+rR9AepuGvSPfcVZohsU6Ti/wMdtC88dv91aX5GxLkGHhy9lVoegYx4NM
Awp4/tt0sBjWfoOOjvw1BYs1kj5DRE/fiMmIYTpSQvJ1Chfe43sMlAQUmtr59QkB
gjXhgRFFcAaTxIqt7dVfMEf1vFNHlj/8jrVfYlxcVO4Qvu24bJJP7mhb3i7xVC/g
Mefwq1en4Jg3OM2pCG3H+55v0Q9OwM0WrwOsZmjEOZbFqvTB7rq7Xq7Xsl3V8jWr
vhl1O8vgxm2EBfXlC1QAb5IfCvkpUhUlvE/pCjsHth/7Kh+wy1wK1Dh0of1jcQsv
0E9M7cINDPHvwvc+2iP8anyOe0dy80etDaRy6OZVFuiXEJ8ARqMHJGbgQ+8Z+s3T
2+xFwAnwj27qDodLRtJUYGIG7Iw7sBfWBklZRDbREa/GFRmLzlknmWZCKQXni5H3
V5niCiXWt23uYL3WhCE/mu8+s8Gt0QrDQ9/+ZP63sUSWEnxKWKqCScww0z+O+diF
NoY1Ww/IVMMI3VpEdpHSBGi/yespg8ousC4TW0ErI92Hv05CKuTcYOniD0IjXqiS
WPfstmVn5IV7FwXZ9uglsswvPUj8YOgdGWEF4VsFO+kI+/3dV0ty4g7gY7/u6JV0
bJS8LAn+05PEq9XxqV9Ec2+9GuqPCjBFUGfB+13q5s0IsZejaslwwTTlsxVfKuOe
CDkOSnHksXF3Z8NZf7bic3GGBaFkM+7rfE8Ykds/czxdKVNji1kQOSBQQsWlRqvy
cfnUUEgy1MXxTP5cnAMDZHsvYRPqSPH85B/aH91cDCtwqJLSX+YEYM31MR6x1cW/
tVC/EXEF7xqpdO86QuMO733iT3r4QeUpKdzr58M9hqMTXc2Rx1lIIysa/pQbaQ/0
mk85Yzn+AHdOdQlPtwkaUYbFhCxpnMErehw2nnXsl05gQ1zOTIpOFZox40DA4xNL
3RhN8Z3wpOM5ParHD4nWcVettIgUiV6JuTinEw766kErjhVwdNHqskpMF/Ln83Kg
/cajAgIlrN6eKmY3/4Q7p//zA5WUGZGfze6APNgb0PQtax3ARZTEoSzlNqmr8v8x
tVeMLBLPN8Ywiph2s4oeUGdVd1i8c0nAcxbjrd0rWWXke1N8IQEYcdFH1DXmgIsl
7qkUCQ4tOFqVRN9g9RyF7yBSl/mHizHbSE99f1Wc9ifaDsLa9rkQ9Q3YMmjq7o6n
z4X4dqseEKdtianjWjhppGsoLao09uHASTeLVGI4L/4wql0kEjWYShDXJjxe/Ri6
Df3eEbrTbb6dd2j5iCwkoJDvNk4mQAg1XlPhmkaPWfFTgE3XtUdF7R/5aZC/6EwP
bm3l3MPbafz+lg3Y7dKnphtYwWYvzgmRPyUFhpIsSQtr/sLZa2r1P06ffrHrtF5M
pimJc0vY0LxV+xH0RhP8kThCS+FeYEEffXgNiDTvw7ryGidNCSdKQS7qq2HJrpwu
31BW4LHClFvTg2eUk7qrldydr25rKhiRgaNUM9jR6fdGAjC9fyl9ep6nujisgEfo
aQ8dDN8gxJ7TRwaK5IVXfIDlTp0RR1pzwawL1Ey+72twsos07JCDykq1oPyn3kKn
lOyansiwB42EUT3+bwPxsBTLbDvnKpywthrGPFkpgQKrWBiQDceFFSTbviHfUlpr
geMfZP7IttQvuFdGAD9R11XbsQLehtdffFWBZsD7PIoiZAwyTDehlnj52ruyfkfr
1y0ZAcXbkB7mCJ5hxi4t1kDKHC5GYGPd6oJlTUR2MM/pDuvYZnhnBgRZ5expiIZC
BOwFu9ghLGNqRQEJPVd9UOZ7Th1aKdVp+Vi45hb1V1QKjXa8u2mXXoNzsKVdPQy9
cMLO0QC/EWQoJi3N0j+rJttNxI2X+579ieq7/QRdRoHS9AkEs8uJHpLMF+7n4gsz
esxf4sLH/m0G7rSMbz9olCR/1SL9Xd4kJMf/DnUt3QY/Z4GtxsvpYRk2KdF1IST0
ocyailQogwP05SCT0PB53KikjpUrpki7P84P9PwDFrNJ47d+76tBth+TwcyNrMvz
H3aX44gjqgNxoIn3T+PY9mzbBoR2QAHSzX41Ai+HBpWpgVsRX/xBi/X7X0IUsE9T
A3/YXkHOBttKpMmIcvdBzvDkHgwMeGOqqOHlmbEr+0cr8/M0yCFe6JIOCseKB9R1
r4TJr3kRTc7LcNFLk9tTmY62LytozVCppIIWdBcaTGwHpy8Kal2a+IiWG0G6Bkln
GQz/CCwnpDbHV7DmrpRljoPm6bx8Zt4oLjSsCQuywYuX5znj+Zw1+6vfhmVVLxI4
kQgDajr2tk7AHEcZoPJmuMmEH4l+F3GNv8arZtC4J2XD5K5VDTuNHNU6ksGDlOou
bmtYF+NBp8wGJzK+c5kGY/SSXNNEzmzGuj+I72lg0o+6xduS2ByZOWB6VwERq8Me
D1szjbUvbboJii9w+1S6UP6pXp7QdzZ7Jgidg1s9WIM=
`pragma protect end_protected
