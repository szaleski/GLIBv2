// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:45 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
YrbcFaLR+repaTsR/1kJwzhvKoDSH8PiuD6WYMsZD7n1VpqsGF0jD7XRUmIcGHmY
DFGU3Ga5JaIF1uXcu1DOkIPXGUt8e/WZyrHm9Ia4rgErkroIPUMl3FffGpqS/NRm
IAVomC64zbQcC3Q4PYmv/F5L7rouT1NGEqCAYs55t6Q=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 9632)
Vg/pR5YIjlnrdMzwMkOzDQDFFbF3mTLNWQBixESTbhkmfF1lAEUreykW98mhLW/D
IvEEGqRnk91uHAhH/QypHnED7i1A9TYJV+v7QLwRmK0XPoYwegByulzrVWdqV2CA
9eIhPzxDL/jxmLRM5aXRAJ8kH/Zk9vvSkD9BvHjM6NA1kIEACqqfDBSPg0QPOG0Z
xPHdFUZFEDlqlQAZg3+28E/p6hvcPO+mjI+J02/u8QcIdOWtRXtfiuu+afymDyJn
57O1S83jnDF0p03A5ZOBRFX/F57Dcv7xmJGo4BF7KjSpK0yFydRMks0t4KBcAjMf
CKJb0qVKqQEC31RMbBbi1HeynPOVn7RA0NNdC4CcZJUMovPKa7L0JuV1mJx2A7yr
bDkDz5k+eIBMPM3P457wZOAoZOKvdtNSktu67QpytMP6fkNXZKRVnbHzudHKoQ5c
uDi1rsTvqAEQzqPw09KhocEiT4fhjyWiZNAbwnMQzTrXzvtdRKzt4f4VN6dNHzUC
u3ZLaJZNYA8HF9R2yw2iiFvcBELCP7AbmocmGEU0xN1xDw3vA4hKkZT5l2kKIt2m
QmYTx0uFILsvwXn5NcDs8VaFIiCMb0RwrnXhsWItgx45wTuVgPw2F44az2tGjeCG
h6yjIoWTfh4IasIqqYnOvUXE5SuauxRZ6yXn8bIKXqJ9M+CdMi9gQ4lk+0yww5Wl
f2K9zxJjXCjN/xpDYkya6xG1I/GVnKiBA8+7Uf0gVnZB3/s0S5fHRoJqV64nk22j
BY6fQ0O5NGnPMy5gj71S6DZN2o2PysknG1fHW8xpjeBvu1YaHDfMu5gFdDreBQye
at0kf2dfVZZJz6cXpYVAUL+IGg298qWFJ+w+NC/aLV770FCx9/ecGiVFz79M41nn
xVf8SQNpalRLbwICGNGhOCAijraqP1tjhi2wjs5j6brUK7D8cn6Fcz+pj7k3Fs5S
iOJAOie+0KlmgSD4AKBh9rCLuJyn8CRCM2wDBRXwagpeXQQvkQh2zE3NkjExdw3D
bwbt0bQXvXhpm1ndbK7GaYzXfRe8JmAJ8lqYSfDyLznVCv+8jgOVbSx/nLijMs+n
ZxQuPFkYTfDriYrfwdx3U9Xk1KP/fhjpXEIoSrkKG2sYIlWCrVSlP4S84MzFXgJ1
cdZBZhS98xed0+qycWEMgCZgUEScGv1yqeRvznvtsGVvPUguMG5peT21C9NIkwO3
2pIpqf6OVwMjNJttz2yf9KOPVb5qYV8Ksur9GWRKyxz3e5iOQ3PR4xg9kmRTjo/K
5Zp0jHBW39JGtux8TveSmvmPqKrM7MltcAhTu02PHpLMOQuQVGa2HfDCB5F6s/ry
/z2l55kdH0kWD46o90KhoSgLRqmHyIoeqy1Ny6pxh5qD53qk8fOA9FwLMERwcxtM
hbKKSa6eohMe/JRI2uMM0/xFQJUBKqfQDv+LfNpaEaAUITWiTBgU85km3Ut7BuS3
SX43MRx81wkDpdP9LMIGYH1oVuKXUmAbUC5nxlXYJyTdPJ9CI5FSSn/16zJ43L5g
uWgpioYciePY0XjWbipT5DYgxa1WyE1QlRpD+DygWJigA6+Xo5Cg7DKnqOq8nUF5
4/idZbPb6bxQrAaHs1kRvEkW02YWiRBdva0ugkq+nxujVCsPpJTeEuV7uam9SV7L
aZhIYhnRmU80knhDgwo91L/o8m4XG/BQsty2GlAAaHHo0aoiO4bWAzEPL/EepGxe
m27/uKmEEnXBbY1ou5ly0kt91OIWnnoIbWOOA0LOCO1FgPJR1EMKYXNBOgoon2mC
1C/uISY/ElyLyvF5h0/wukIeTdf44Ex7IT6WeHRokRHa4NG1cCbtlwT6XfrRXtjB
qE3t74k8gN0OQUzqwbJ6V+9PBKKOPqtgirB4DVDhUnX1pCxuMf5aC6h9mqH/TYBQ
Q2MPB32ZHMOgQRIKjGTIJ0326pn91Muf47zho7UwsvtNsUagDejD9meJlVBwHdjL
1oDNXQQG2RkLHV1Vnkn3JCUBKzXMTLkPZCsIb2O4mxzykuWAJzTpoQpWm/pQTqtu
OzAJFwmIuqs1BWszc/wHiUNPJVxclb2TczxAa4S6NrKe1BCFbj09UKIGIhUptufV
x20mMochV+6HNLdmcqDJVCKVs7L2+NwcnVZXCwSxrzZ7/BSwpicXtLuQzR0/Qn3X
Nh2KCJ7hOrmz0Z0pQaEI5kAUz5K2U/jUNiKBPX1+OFI1JXsKfcWLyaAW+iaPxFYi
gleTRM2TeEX07+lwO4W8nmwmxjPf1nHmlbleGsgsxqX+okqlf6598cbOP+T2i7zZ
4abgXdXIsT6ul5lhyaczH8CpLDU9vldxnXf9DW3wZJQgT32NFnvpMDlaZImqonM4
8cE0LzsfsApeJYfz3fJtsw9vO+08GRPzUvyfioHnGy2zzv0F6WiVS1oqgIHQ0dY9
b10vD9TXwNF+9aPKhN/f4+JLB8qehvS9P/AOME4HmCuRu04//tuOgAh9I7SlxDyT
9Os1hZbZy1MwyPjkc7TT2uBtQNlUdoxZ9jlMHwVCvcLCi4U78LLsFvImfI4QG2/H
jm7ZfsiYVsVhZZkSjJ/dfqA57anDTFu7h8QO9RSZDThIDjSn+kqLeWcqLRgUfi6o
DEKbX+sBwa3Fe0491NrwTT3u26hoJ6AjrvZ10r3Ho3zMCYiiWGIhhJ+vox6HoUM/
p+PKISwL6UA3JyN2+nljkU1EzKShxQ6qxpZ3V55zXh2KaoMyPJWMvvDpvbe3tQn+
6OiMIn4LDwkn8GG7btl3Lpj92GhZo0qx1YHB+vaeCrKdAsisacmGkgPjTbPyjbU9
haf3XkCEng2Be/qg2LqgWQBxvnrGzK+Z964+XctQm0N1v9Am65VL6kQ5QAd+aYpp
wR/CokBs5K3NjuJJR220HILjXAVfwmeZfvnFtdsGXJYtBegX/mFVkiTu2NBi8Vkd
5MI8GtccEjUlZDBKUT/ECuI1aYFKDjB0pZysoDgWLVFaeRC+SkkYqvWth2XUEM7G
WVKoRRiu+oJ0Kz6Jg2seZfGm21NQPMjq5hfpdAmi8UyGZnnEx2XUQ60BhuX6iCwr
O+qGw5lkE+Embnk49BGQHrw8au5TiMWY0rVFKVkyjDHDWHjszZqn9brvML4Po5MA
R39PC1RXndEQzLG207rnhRdTjgVJCvVOEXsiW3Ila6iOb+iVLEywqnwaHU8Iz/yj
kfIQGoatD/qEDkXxQUmEAdGtRr8cvfF2w3du8f3ydfQ+OKjorbzPdrr82qgA+FFm
ZEa5CeGBh31hfmmHHdxocZbILOHNs0svbW7okizl+PvQNUmG77/JgWq9Wa/iBaBp
dUWa9JQJb4YOP6DHQK6QaNgCoXMVpw5ev9l6W/Rjpjxl2Mpio4+mGnVJe/uuPggQ
57qgnRVvGsaSxzKETqlsjWQ7Fe7/H/LUYjmXn92nKV6t8D/K8ix2bGvlRinerNhK
l+AqrwJGt1z1vxCSMWz7j2tikeuoab9ck3T/mL8HZ//u8ehnmlcGbIacrO1M11UP
Zc4jC7IkLV2/1rtI8f/tf9ZEwtT6gGavJyQ2vKDOe92spKL+Rp+INlnQ6g7cmjGa
Z1yMIdPlAaaqWCq7pNUSPoEEVbiBWsmowLIOpoLsKxtiuhMGyuWXAUxE7WIxxAxQ
kclVj8VhVcynYB1PT+IvKYgQSLHz6JYlPEjtsQlrpLiYNsRmc+QIFnQcW9WzShxp
wc1M4MqnbVnXvVGU5yQ8TMOikuKOoejPNu+RJJlylHP+1+o4ielhMy6mKx3hEBZQ
NzVLRGHsG0ASLDhERtWv41oWJ2GE9K+K3cSh4UQL37nY+Mld14TUCeKkTEFN0k14
hqZ4NbUBVbOKHWS0AbvpbmDDZd4B936GYG5q7Wp7HagvJDHl57Ye560K98b7ulBQ
Y0cbn5mbUXUlEkHWEDTHXMUmp1b5NzJRV6DIrQBF+oDtfyuYN7H9JWdPWtaZiyx4
dMPh9zn0SQwNiiDoR0JeNSUemJ3F/Xf1QZLCKqd81aYUyIzpu91SGFpgb/1+umsm
042VyzVyFwTi4J6+MB7AiNPtgKTfSh6xk1u++HCKu8DhS5qPXopy5XUCQOaPvsED
IvUmTmTv8G4kyRG7nLfh8jDfbtEGu2dpaelnU0aPU0W0QntgNVsJzKfHdHp/vHsl
N1w0ty2QXnQ++tnRltYyXMujiKveNlafcHVm/qnglIPs18heU8AvU+xIzjSP5Jck
1zdoGeQo/06bqot6XZOA+DLMzbd8A4mn19FOuCrhQpiKmH6ZX3srE9IoG7FBn1fp
uDCKjw9r3bmgNywsXP/YV/yNsLmeV2udxGn2YIlywYjnnG84+b7Fo0bAVN1QfiA6
bqPmuIe8J5wgI6E3+Xtf9y1kWjH5tMeDzaV9wyCt30mS8Z6Ly2J/Kpm/Hp+Cfr4z
9HfUOMzdDPkqXqEKK7yJCfCUi0cQ0KxuMWmqNKVOgZHYj0RTcdPKfqrod5A/Dqnh
CFj+8SAqB6vBIlxDf5c5vfaSRgihMln5j8gOY6IIm/3WS7akjD0m03N1FM9x1j0d
p05czy2o0U936Xijhp/EUcWvr7fwZ5Y+yy0ycL5RImiUrkUy1bDfIvVKOB637YXV
HQTZuCxfZzde57KZO4usprB0EyY0z93lF4dCVAvZXxG5fcMcnQsXlWQU/1fxTW4p
ANeGXwzLXVlEXrgqB1huIDAqHgpUBNIU6xXDIIWBcrx9x3FifEHUhi6Jq6IaOC0m
78GlRRuU/DWEMA1zY+GUEvhlhdXQGtohqNVwU8fCgYjxp50O0BJXcXRQ+PmDoiEe
HG0Cc2lGa5kWSMAY3lVTaETc+fP9ytmL4leddyW6zL96dZ2JKVN45XaVFNIsZfFB
k6ftkG9WRtX2ZLB+I7mWDu5uozqAM+z1C5QYBekrb6lk5WrBQuZC6L6D8GUe31QG
IsBvAiQlEf6j6vBle9IL7Mm1lbXJOPZ+gPENLefj5dn48clJl8mJz4R2xbMmB75/
4+WCfj9RN+fI+y6xvcEfr0eUi3J7axdJkD1GKC5gIRUCWnn6iK6I79lfwNnvjTX7
0c2CahQL+nuHV9Gk4Vjk/v4yEi1EiU5uUzfkViIx/yzeoZvqbgGHDSeFGlAnhxvQ
3oj6mFmFiDuU+O5Q180Ep0BBHAfEwqF7hD/7H5V3pahjNKtXPJnaCo30e2CUc1ku
vatNZNcS4z+3doxLx42Vyvde82CnNukNZKKZqCm3IOFXM5Bl0fV9eQyLPmF0kpud
ojCNkQ3VkRa27esMAygGjesaYxFUdAqDKNksOJCvfvWKBjUgdX66NbpBRhJcEuEP
iZ49/4ZGvB+aGA3hWc6mC1zmE+rMsVVRfXHBezXBn9ECu+bYOBVUKgz+amOBatBz
hgZOnHRKwc699Cw5eTOahJ7YvpOz4XY5Pwa+dFSqupFJcPzXBkMtDcEa4MMiwGx4
7XBt/w0eZthPd+8kxm0dXnOOfszTFVvgzj0cQFatOTm4ZxN562kEa1qXA0UYf3xm
LvpTenJqgeaof31X/u/UrzkyowW3814dEZ8iTayrojY3fbYCp/vi+Irbl4jY7hZ4
UIMWllNzgdJHRc8Kn3ozIRFfJ8DAAAxlurKcmgJovqG7g186UsyebUOjr3TlpcXo
G0n3sj7FKdwNysj6SacEgrNlgQWTXaiyaZW6ZHLPR52SAEvHNysIUH4BcMxX7Qse
VTGgCzAWhpQkW5mbVQxe3cMJjGMZPUC22m9Ix2IJ0K8PKsx81InqHdQxa2iTSBcU
WLkjJcYw8FuhXCRkuNj3nt0L3B/26KhmRx85jrrECN5unXeKTWI5bsdDkfiHLWLm
Ozp6Yw1EE768oOve8mjNhikstCL13mg/cBJV8+Yfn9YbjteEhhsGv1tJtZIKIhA8
6athos+AryB5GB4tV9KtBDQzl+ZFwBs3CENcBJPANNHXRuxlTd/Z3w4eZbjFu2Mg
KNBWGR7BRoJ0z4BxmSEXZrv4E2+s0N36v4e+mXX7llrt0Qffz+Cu7WghlYqr7wAL
r3UAOSfFLuec9zDxOI89901eyizvTiqQwvkTTed2F67TAvaliUYBRvLetIglMi6W
4VeQz8qw7ro/Ugs3xvQUzyp2tKSpX9JR1VF35wIcJb+63hccXSMNr1g/ljEhFiGp
VxBKScf1XI8QtVtuk0aJeyRuaXdByn8qs15wxAVE1GvcZmSI27QN70SvM5p8SrKu
RmX7NOH6S7UhfvJjxKYHMZJhkcqOwNLXK0zmMXzHiTTWe01xLzr3pn5t1un6E/vt
yzIC4KetmOcqB+D8K370CGOEUKHCO/cDBiGwaKh3GNuosFPlGsG4JGUqb8qCngRB
wYn2PysdlxaTvQHMHcGGVTAlz0CqGgFmbBMbukM9ydCDNAz6dw/Y9xagJjOJRlCz
Ws+o+VTkAWmi0ZyCrEhCnwZgVqVN5oOUNJ4x3It002mDUZaisKkqJtLhD4ej2VlM
z/lle9sf1bo0DZ72lXIMMvz7+P2vSPOFt6qPNB9LddNyqa5q4ab8ow7O8LfqG0m1
dLLq8AE1DoHAOVMXWOR6qd3l60I51Uif9NZw3OziFV9qIWE8fQZ0Xw1uMhukNdkm
IoZUQtO0EiSa7JiRGfF/BthX/CeOgvT1GJblQa14GgmhS2oQ23rpdg7BPyQCety4
Vip0wtIUNlfathFkeWVSO8U7O0nFe20szAeXQwVy13VwOt3YuKZ7kDqtf3tjDoUS
6Zly2I4XsBWBH3RJ/bwl/KRwBHPxhKBIvkCpd6AuIDj6ZJX1VPvVlXDYURuYQO0j
3zvgfo/6gqUcEi9ktrr0bt3U8rH2lUiQX44yfrkdqxRnUyLwAk5AxHBVFyqDMyQh
7FslD8Zk++uvFHM1LBndddWNU9313Ry7/JcEo9Ko8Ox/jZ750k3DOdHXQGDGSY8L
kQRGBSrGuZbvh+TGcdZZSAMfc01WUGv8BJXDVsIveCrDBTx1o2HxGztN651kDngb
agAz2UFGJaEuRYP5+az4lpJrAl05btfw9e1U+b+b8D6CrJUuKRprdMOTtqyFUcRQ
oRAEySu9I7R0+4CoegEHe+UXTP52l8FQ8I59OyHWvWaQHJ/MsM7eQfP45hO9bcm/
4zVECBydXPNXjq6E4u37lAaXYVnm+E5cUgAVWJgRXqXAyzTwRuN9SL4kgc+aUBxl
HmbH+5gCQ3r7mMx8CFSIBlO1IqG663Qn/F2JU/XunVcN4XhnVT3/UIpZvessGw4a
FvswAM1hPsGG1Xh3XdWX8Lujgo4vzG+777TJQ2o6jFK/EYteeW6stjSHRhwH/Uql
nWP/oWYU7XHqGNxBEOWRjlcTR4Q+oyVtn8/Kass4+r31+2QCkorwqdnok1WG0lgs
6YErPVjbmRxOw9tXcN1GNY1EN3+3TfHOxU/b9x8Cvu05zigX3E7VIISnoL/yJNIR
WfCaDpVDMcjK4aCtwGDWiBUxvb/PI6ITgOTZrRUMvHtUwYUHGdx17+Z3MNx1e3k7
bvnq4hHcSb534KAKFSzFQ4glYKsHScQbmC5gC89MV0oDxZoP58/+khvq+xJkY3T0
rVcK2IMC34g0Bli2Hl3npC1UHoS/ErDRItphcGYV+wKilizPm9/9if2squwaqyPy
IwyFbqFDr8ZQgCvU8c8eCm6yheYsXAlH+ujCLysQivYIneisl8NS/m8qODf6Zq+Z
c0satpZ58oA7/0OmQG98aJuRw6hu5UhJk0JwYjim4RuIlR0ypO6DsiRSRjKihiCK
bSPQ04f2+s5xEqJ8e//GnnXUdIoD+Sc0ZwPkf7+nsgMXPIk09r8LIqgXAg9xnPeI
QaUsCkW1fRoPi6QLnmqVqrtlCJ1b9uHfAa/7P2/dEaWtkWzLA7lm9/wz6BRKmnme
JcJL6FWdW0EwDqKAecDAvdiNOE5+LvwYAIbTmLC2fhF3bPLXmSWmbyKn9+aOOtVa
snLZfm/rdgvqk7RgZ9GmEMMjo8p8lfqI3hzTKig4O0EuVHmAL1VR1nA0hjAqZq/0
R0vaFDHiMRh72NYqZGKpfHkkMoQawmB9E81tVdMjjUGzmSKvPD9mBuUyr77m940j
FiMPi51B8yU+8HUW8sKFOyAB8QKw9yGBT3iRlrX0cr28DkBtLqrfoYfYC0Z1x3y1
Du8PpC3ZcLfPvArucfb+lUF/f2vlkWOYqwIODODb6DYSeV60jcB3B3F8ortTcu1h
VR+/X6JcZ5zjZ9Y9qwbPEn/fNyr8L9FPVv9ecUKXvGxFpoYfk+ABZd40Rzx0rZjE
oNYpbYUoJsK3f29EkVzNiGnmC9WV7Y+q2hkAv74knQwtzP6jsIsCuyYWTkPaZava
leuqryeA/RRDIHscipkSe3yQtHzb5dU8zG74f1Kqg43DoREbZnb1QFV86zz0odUq
t136d9hrJj7kZTT9cQ1KWYGQGpxImAuHmw/NNkr2YONWfZpX6bQtgLJvMu3Hkt+t
brbpFxsnH4NADaqPgoHERcLLY5/OnfCLEKAj6IDIW9NBJ8mqI/DNvzCaNYdtOAhA
sjvPIFVlG76SMx0oVS4/m0MT4ozM23VlML4ogYOA4nNwtbaEmIT00Vwa3k3ftft9
n8lTjSuWGEljUnl2hSwmDPS9bfZSZtTocHPmp0cP9i6l9HXcSb3H2ftfeo2Qdw2D
YX7XrTEZi8sLe7Oi/Bw5qzUmzkC8su8nhsMo3nJN3v5EKOAi2FlvmndciiOF+v5E
O4FAZIQOpccgAhiTmVfOSk08Au3WRqgc+O9cnJFvRKHBrVzQR8HIZ/oKy663HZbo
w7RiqXjD42SfxCFNE2XxaaGuKXB9vpstnrm0wTZgY8OcZS59n9ucz5J0U07d5R/f
48SNMPb1S7yurz7SF6d9tpXMzZDcQTVisyvq8C3zV344pffU+6mSihPzY4kG8czG
pcM22OVc3PS/xvRGw5iZqdW21ck9CtzgEKlNItlrH5NWxQPF/+bYGrqst1h9T3N8
V9XnmZgnBLp7BAdqXD3z3BTFWb0kzS2cHWCNaTYqXN4v6JiSuv5C/lTG3jfULtW+
j+mj8KnSv+JoC9XIXDYTME4goa/sk4Tq0I2TKC45uvYGD/j9j/NovkYkbjgjzvP/
y9fHhA/F8W+eY0ukXMzAAxUy5i/L3MfbLBwANAetDM2LSqn/bC46rcIvM/YB93hg
TDpV3ge6qbOBGzSOWz4v0FS6om/COLrqpQujbMq9W3+GZXg31ANAfU+rpnVbllXG
MiAn47Z1BDmQIZjigCVr9MFKJ8G3Ln09GoJS/plE+TLyaA0M/h4br8kFJYGiNwG0
xs6W6qtQ7YHQPdwbCteYUUlhbdqksVBN8B7cbR7OD8ynL3sGcXWmDeH7q5/e2PAS
ZD4OuOpXMzHZraKYbCxfUo5O4mdiTNjdQDx2sWfrpvAtOMZJ6JU7p+4UxnlGu3Oi
uq4JqmOCy9J59btDVF91x45CqkLDGx5yWp0eQiVhgpNOmLjRoAmQYmJj0e2q+/K8
eg5gb8PL8mSQ5b3B03zJnz2+LjM1VXHDGJXilsu2wAB27T66h3jpSP3NL2MOj1Jq
vKRQwGtGg8F6Y5VRnweauCQ8RSG5Dit8OmGERjqcaNMprd3cW1HjkDB63p4E2Vpi
Xzmxs5kzxO38OrfAxj0IUr11Oy0Lx/Itb3Mq/cdTpeCWJT4tiRJN4bLK+cAw3okl
RjxmUL01zs5O/QHETtyPHbvp6gVlGL2fbKvOoNYKteZ23/h+9dWBkKeNI6rlLqlR
ld93LQ3tkGo07hbZXWI1JiWU5xPqMUABACyTNjrLD2B0ADVve3liL07UdtHcQlNv
6046ZJXqXcUHXnTxSEUEjVGlSi3iR1OJmnnzPocGISfIWws2iuelsDH6rNRYfEjR
0RIVej4uFS7EcfG+GLO2ToVB2ei2SEgJ40ka8JgEmL5mqZLRrPpTBIFqEUoBznYN
8k2PrB6OFweqd5oTRmBj2hlf0jvMoaLx8YnlHIoWRyuZ3lA2TBpA7krV0Gsj/hlV
G4fo2YbuK7FFwa2lxXp0H57zrRiBEeisxPkLbfG6ZRmELD7LZHZG/jorR8YDqLFr
1Jd6eTdHysL5gVm6Rmbtbl1lJOsJ4zZ6ALFSHtx3V1arH8qNzypxfrnXiY/hy2Dz
4zcUPvCwQHdNuhUFplRwLeMO0jl23SQjzLWtqaEww8bsFWc2mQ7tdOji7DJMTs2K
TSKLOT7kINDWWzTTCy8OX5yH2kasK2AYlRVz1I0b+KQBwJYaOOMgi+5AWv1Yna9u
jQTNeY5eh97Wk+L2L1IUy1HURSaKmVcnGACz9WQFX1HbpQOLi961V05yy2M8HwRs
a5n+M8mOOdat+UZSTO3pzhn6Brt7M9epJ1iRBg8f/tNyjctrc5D4nQQSCcuT74sc
2HAoTcD5ZGk4fs4ND6aa9yw13POZHiqAxSolkDAvcnv18EN2MV3JoVa26FG9px1b
f6BUeIjVt4U4PkfCApKkLrO9IMd56LKJjvy0/BFUjKMnO1w/yS2nGzRkB3nMTQix
kzZHi804lcqTz/zRjZRXI5jkqLPE1HqGC6PZUV9Jcj0pyeENrCSOU156aiZRZLKE
93nJJKsDbbuyOSts+Ws9Xx/Ofl4EinAcTygwwOz6j0IJL2I0JJahVGMGiJ+9rr9S
VWoRE/8/zfFyNeDNcLFAnpTy0cYxNyqV8D8gHt1mqmil8CgBgziRxOWkgdFj4uhZ
b6LGNtb15zAgEuGS5IuftHOrL22vUDN7eGppbcYw1cmQ3hHeIew4z0gZa+RC22xl
qlFL77h8Jso+BCbbrevjx5EHwSh2PJkili0s2Jtb83Y0l1vEcKxIgxb9pM0cR04b
oEsYEYu86iDXFkZLHe0mmQPn9M/rPVc9+EXfKkcVYLpnx/S5ZxLUlvque1lGLtNO
Y+ZPyx+YJEMB4wra7x0GhTPUneiPyJsKr8VYpmScupqZNIXsn3G0n3NC01yWF5e1
+ovcbuqi3yQ/oH72dsWqkig/PZov0gcxjq5YWGIaPll664RoR6Jxwxac4vYNRjma
X1IKKNpx986bdDqLZLav/NOab8a2OkrldhsFoDGMyVxYkhEtsH+jD5Al18FB5r3U
f+lmi+f7Jhzy+0uzNztO4PRfDXIT8b4iwKTNNxmaq2AFp3sP4r32itEUc6PKfs4P
06FZDzlNRa2KUzdLG5vAYdiVUj+4cJkNvohctLKbBuXuoqtNOP2k+VoFOzfDcYmc
jUhDk3DpZlWPzMP5jtVTmz16OZ+fYSzNoqzFuQiiJUbr6XMJ0wKeWOSlczFkYiko
iVhgxnNBMQ4VJgnHlcjv4MHWjEObG3E3hDbue3ytpL3YwINbNaps7WdAwEA84AxV
+KK11GtrNFIrAOnCEHZMbRNyjjAyPINGucAzknbawmeUNMMgHD6dwBa/GmWtenwb
hAcX4YiBsE/h615dPDtOi0XuW5uyEuURTIIYCZzkQmpVyhn83VgW1TKkDiDVbQvV
7jTeo8JQOV1LjmIHLqAR/Cnb1xtw+4mK3Z5Sn2A9E+W01kFq+FigOuFV0N1hagf+
K2MNXE7e9enxCYO1ac++2Oeizpdj4TbDSIv7n0AhZzNsajofz+MN0D0DGIMXSQa1
j4IORBQ7+8YawB+2gg5Jc7pMr2b2PG2Apo/lwtaOuwC1ZIMKdQRB3srQpQQWMS45
Qr/lL5XQWxqCeKUgSmhXD/FiSJ532DQPDIhPML9zizxlu3x9jEsZOD5r8MYfDfS9
+3vtOyfpVI1cvlLM/Ocu7LHbRZuittWZCbNC0ebjVXtIZMtuQRLuF//N5ibc/llV
7B5WidV0ufop4v6GCS1A2R+BGYhUW9Te5eAcZiqjDsypdEqsjcfd/Si1yogXaUmM
14mR4s4QXl/4evi5Xm738xsF5hs6z1qn2xRLk/TwC39GUvEeP4N++tnIlLV3/xof
K3BQEja626nnwfDeI15V1unsPSC6bROHrU2cSB1aCkXE47LK91eyGJYLBxbceCSi
jmg3A1co+e7yVO90GS2/O1nfFkbPC8Q8ZylEJCnXOsM6CMlPmyhd9XZxUE2wnkWB
gZq2sF1+MK85438FXqX4GQdXj/3Qg8ebnTaOll8kSbXTf8d2i0w0tIJYZz9rKbJv
E7DmqTzlrMLD571WD8Vgpk/x7f9z5hML4EDgFQs7oKBrRJt1hZHo70tjBfcapJrb
8XMRFnl2aaz47618UYfA0hQCDWihIXoweWjegojgmKUz/ldiyQbd0I+ZsGlmHNrT
vNgZAIQYxc9pSyI51Tq7e8ik4C6mpGd0W6+eOkyMxPwH1CXQy1KJKzsJT4zK2V/e
XoEfwgV9QFtDIk3wBBKidwt2DB+OEl0v8keg8cIHeMuM98nhuU/WDcUseW8LzKXZ
dGsAb1WMUpN3OPeZH/TF7uJO72cVRFJwph9TOCXhmYZSXIOouNF1g4QsT7rOUs1O
BPQeHFjv7ER4EN8aZgH4h9j0cZBEpeW1T24o2MYc4Zq/iGdNul3XYdcWn1FuWHZ6
s/6MgPeULuQ/nI0Ye0G++BR3Xo6NO1/n24FaBShuwBMBsSDtQTGtgHguN9NsoQtn
Okv790y6VjK35LuvUwSMOumPecD7A4K3mSEiTnXTojx9yM+hKdRWeG1QQDwvlj1G
3Pk04cNLqmC718Eb3tPWcVaorXiiVDF4ezKakjIpVQ7hgIjib+JypwrC0cu7oIBI
JDhKT7EGCp0e2WcCKK8BjMtDQYdPouvnOEDHWlX1DMbMtDYzfyU1X5G2hhiWhBPr
nz8r81lugBIA7MrwsUAf1VlHUZSyUg5getYi7KM9XTNi+ndP4w+AYpvP1bbquvDv
qWkwQg9jSkYuj87tj6e9rDpDs+wNeEXLEFug8v17s3M=
`pragma protect end_protected
