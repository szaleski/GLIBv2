// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:52 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
D4w6r1RInY5PdBmKDF4egoahiz4Z8ndan62qAjiKqSngUMhEqvjhYBfCHz9BSQY7
id60Cf0b/il1JNoOtC9nmAB7csZ+7ymhp2WN/zu/wIx4Y/paBWJw+zTH1BncF4E4
Xo+lga/OE05wTIAc8iaxoywf8W2vFO97jHOab2UgMSY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 9216)
OhOx3TFXstM4YzdQ+j3LOs3OoBAogfefUf7tPM6LInxf2+mgDSxvCuxSUOd3VGEg
KAlyc6mtVzbx1YyY7fRM/krKDhNA3AsTsVXAvqQw811EPOh9D2Q+PPGy1jPIv9oL
PE8NYDcP2cRPGWyCiO9Nz1XMIqQZbQLYBvvXA50yo7eGlcEKzRf3pbt3NjVuBVaQ
TjvgkpJN4/w3luBOd0/SNlCImCjQ6Q45mAYvFV+rsgyi/R1t8kqRkyQOEjEHsDrN
Ye1o6ZGwz1TJuCMr/schh6zrGnXm8a8GV4QJonNUVED/08LqSDkyc9Euz7SOnYh4
ARmgR+hCwFjGHkxwmuZcjnFtNI5ZCnSs/mE9+qm75CcqNW31VeSHmgP78FOgbSoj
VIAttzaXC2zlsy4PamM5sFmegTRN/OWtA+wmFHyX9JODPh3NVtwKi7dYALYuLCY7
PGBD8+dV9jecaepch6VnFIuTMoV05jyY5K5Jw46+OtFTP2UYVLuWj8Mrj7d9JeRz
gcmjVqkEwbfzOWgCOi+B4vfUhw2EH0+GHQp6wf1aBv1T/hR2J1BsLDy4+To8iynQ
yImNy4KqTkgcFnbYPKCEifU8LJwP1HfH3RbOgCcCWyG+tEw+SgzUNrlVPbb6ymeK
Sn+/gZTVbgw6KZCAzkHw0+N97fiA7c3qxzgd/ZTkl79tD/UAOvQ1T1mAjg3IU1Hw
V9HCF8NY2pr0vUazhsf9ZxdsBh7+CcyK8ceJ9Ykm65PduHp1cC21X0KSz9OCi9/5
WSfgE17arj49IWA/tPrFUuD5WsmDerUDhCD9NyafyTpJ1C9f0gr/DMO0Mqtj+MAO
nBQebNANByni9HsXLHjAA3mN6ZpDJfYO4xUVnUG8xMpI29FuTDA8fgmEtAlTlqED
h9Wj8TrC4Sne/yIGkhhxk9cIX5Cn/Md7d9jk+eY4nAHhKi6DlaNRmBNEQRxGrLTk
jGY5XrXPTAHr+S2GnTFUwFC3jvFGcDLjQJxgyUThk3lR8IjQjOupD0TKNpHihn5n
kS+HFDEjxuODD1w9jl0fqKBT6dzHVcaimj24ehscEFYeaGvLk3cGImYwcqbUEKWx
1b1ebL+3H825tg1HtbUSnrI/Gzoc++qa8mtrO7vRbo9JkJIEgI6fd0MEhEkvQynf
DgtSUM5/SkY8OlXTPsxv7Tp+tPRsnVMPwfdzV0OBCjQGlG8SUk7gtCe8SMw+mEvh
FxYQZaTmxNea7xQ8LnR7hYm5Du4SJ6zwlBD/HdWn2RYepbYL8B8rWcADmdoeKY8P
aI3eHF+4CcfF05K+QRukO7lIsOnV82Q45CCfVAGHts6GLHrftwLdFk4cfzGJtrdE
0viC17pARXtxrp0I3FkU3vPnoVu3Gb4aWOELel9trA9vXvfZnNtKaSU9dzwNboRM
duWNIYbdMCK7egHP+LJrjkCqvqwwjt5L0dBhCeJZPKl5IcjKPkD2lhAWWjD8Yogv
Hwirs0L7+EArDMQ2yTe+5ENSgefauoFuExE3NXmuCUM9Z5vTnQOEtuw69DFTP4gA
p9562rxnmfzKXmYrLBjoSZ3GIiebyZIOWzZ319hT518tjJs2rU2lDxfO2PVH2omM
h/dEmK7v2wcDaWEdm0KwcY/28onQC1YBExsfIFN5uEdpz1tjEV8scZjWWBTYifY3
Ermtf96XTAKE+RvUGnrMW740k0xVXk3qJN6oSfEZOMal/1TBwjCLmHC2O1RuHPEg
9uRINS/iah6XPAJsg1Lwxclo83lC/Mj2NRMeEYkAWHH2uSbO0Zqxi25un1xs4eVL
sUUHuuv28xysguJhEyoHlhF66KzZKmDAUsVf+yzTyp88iL9qQsXzORJQYBCG//+C
zdTOKQOBxfeucdQTCegXq2uAmYE5OardU7+qab5F1ou9yfqZKrapTzrdpcNDPyTq
96eKUe3aSMkN1AsuarXAYKUAr3sjOdkUuYb66/WKkENkRbTjRqY013TnBOepI+6/
/C0uRIJVktAtcHn41ED+i/rq20+jHaOyqVf/eNcEsGslHWt7WdQgg1o8beKpJizW
SjauMRxkKPgGLhaH0a8GicCqdLx/kSW49g6Z2IKhodopU5V8r2OMdhx9WAXYXhNQ
pNdZucWovBFPCG4cngxf1FlPdpiJyFvkTp7aADnPiYBl/p5LrN7mRq+G5sovjfCf
7LJaUO8PX7QjGuqf2oY+grMj3ow3y7Ejv+6tCBA+pYWDWToIrZuT3yju2w65hqPf
RET7Fw8R0NFI4JL7PYgJmxPe9iJmJ0moeOR7fnRVuPl3OPrBxO0akrZpvy/OYu7W
LSnCQ3k3gUQwVmEbyVD2EwzODQlFFDVx+VlPDhAcjQVkjjJ2KgaK1tqj1Y7yFACr
w2iA926zGNwELOs+yfmh/oWK7nBjvIPM4MP5HdjukUUQ6kNtvv3rdT+fe1PCSoT/
AgxBV90msUw+3gI9lNR4ai2uRCFEt4ParXt+7rO0sC26ICTN/eekMqXg4AFI9DnF
uf9T1AoPG6s48px9Yg4gXRNa7BerOxKGBNwhWQm5BvkRjpAjZnwOz7ZHVUaYkzZg
LDVtk46vsXKXARYS+7U9mJrRIV4Pt1tIiX4B2ff32yXCR6Hvnk36gM6XdroZFwE+
mjmYQTghBTEcfijhgPBh8fMXfd5nWlQGvUJRslON5HMkl0FCmozvOZKAU7vCFtRz
IKpqZAqsNVWcnIf/+5SxLKnibfxA601O9NkpZ9EZlkLSXjrHToN1Pt+sZjynpGPm
kElhbA6G2/iybzUwQOD0gy05MN5J7fr3KHzZCRGEltxDy8M5rU22xfZ39FSK1WV8
u35K9wZm1ZJcjCVCHZqti4xeAhQWM2wwi/En7z+auvbvMhQDN9hd29gofiJC5ajT
bG021Su30cPcgvI/ZNrBpyR/8ssFbtGVKhwR7iuoxdYsB5PjmvjqywX5HTqpX6oO
BaBLgsAsvyCY3XJSLDRGy/T4OiPdZumjeeDFhKlvR9YrELKxjT90zOBYY5VmvT0+
Yy/sSJyMlIUGLbNJrq6RTr2UWOMFEzQh6XSAZFlPStwaBP1jdqoxEusfgr6xKoB4
GZe7ubXqwsY+7yaml5T/FVte8BWr3Ml7Ao7MNmL8ZDogsCruwpUdNmpm1UoHlEuR
3WmJEigVNnLm/GWJK6DmIaEVaIFFc4DbUoysBE99ODDPvbxuLDGFLqp1QB1jh1A0
sX5XMDjMk0pgGJxwb+Sl9k1zzCGFEBfNGjG5ePdea0jzW0OPLEiHJWbC/kTqIEd6
BDs0FXOJfTNCGlIQlbML2Rd0sr3lu+jz7XxQaT3lzFiieoFs3UN++H88gmCbuQoi
9cxGviV0RlKLkK4882YxS5gql0PfYJTQR65fz0vfarVM1p50rZMEh1jdSvXZdnhu
Y7/eMsAhsixXGCxrzSX2SYoyyOmpWRCn4MUgvWIwStOgu6Hl4Jysn4C3uQoCLg3U
qwiVxZLmbfd8+mPwsAE3Dxv/rQwYChAdO9s31vbMp0HtFCSPPgm8Yo2UHac7apE/
JlVrIml4rMaSDOtMoOzCwzzv7DHASCp27juHz1n1Hc32CJ4qSTdv51bFkOly/uUC
hJgz/DYlE1VJ+bG69FcvLSqBXDj13fzHepypsO1KaiQUdx8dWVUh9QGl75aTZc4p
qnEF6tr0Q+CA+YLGepUI1w94tYccbZknaykO4thW+rNQwsTmxODz2HzpfaVR5dyL
d4PDVVVJXXW3rFv/EAVX8IVAxD3pp+KxXCYJ0TLnA+CtDAcX9LAdxNRW0qKqGws4
gwoXw+NCvCie7XQRy5dTu7iP2vg6KsaZn+GHKqz2qp034hBPyo++6K5BabOTl812
sP3pBkK+JoiqpK3EMXSFVoLcRK9I67Asl0dgjrmUZYEWcIhVNQmc1q3y61+f0QiU
f5E59bcx7Yj6XMmfO+SW8KFSKLruQm2C3ujV+6IJIQdx1WvgP+xd+SG3QZouv2bY
kiZsNfC7iDfN/vKi6vG8AF8hz2se+2FFcGh0TLPkwkMUkPCka0DXfZU+lBEYNc15
UjOjloBxYBONm4wQkGK93rUFeSw6yfxhP3zbHD1KXC1vvQ6l6n9d8CfW0Q37GRKH
ZIVIGScCbAX76eohsnG6y2R+3VsWJsheK9U6vhqR+r8nRevCQ+oQKPE7wE67N6Rq
T5R2Rp+371RlJvHrCYkMAx51ceIES82sUblfOdZ0o7Z6AlGIW7HgNqzmsQXTeO4/
Hwrg8MXtwEnyquMesYrJ7w9zLTexJ5mpQoEHJLFZ+OZLvTaIp2IwxkPxdxY0vOpG
d2yXkGEgt529CoVz2UKW4XWAPo2sXhITfC+8HA1MqlKVUIJRoxqRk5bdWxtfmvAx
MoeaonNpLocj/9hKNuXFgFAJHSWWqwK8TnplHQ0TUBBBOaU6h5bfEF64CS0kd+8W
L3OhSuHf+IVeviKAQdlXkJgNXwZGoV5JaEaQWQIO1wpD0u+NOhP1wZ+EPtkCly5Z
KjA8rV9PUXemb69f5Kg+xXMFVxBIO5V62tZTHoVcAtJwYfu456hdFyIeDkKc4STz
YxNvR+uRBW5O2W/YsiWdS4L/g3fM8QEJM/qijw5IeaMGVpL3nLRwYpcL2uSfvrvJ
oi0Wd9bDi8lh0Bp1sHkXc4lhT6kUhKJr/nZhj1oYzTwbGobIIW3hIXi1SebfRGJp
g26mr5OEaag4rbZ6f4dhY/NljhAY5fsrarlOOTa7buYk3h1dWcofFrbw+6zDZKRd
qNGj5qmuytYfLaN8Y/VwD+ds71fA2+f5+9eXZqW1yt8H+cAcpBaEjMBkCiGw0vCl
pC5z4/i7R13qj5HL9fzBT46coU+xtGsNjTMBAv5n2BYRQnTseQCVF0bBO34XBTGa
EvB/QaHxTUhPaW9AplnRcq3pwdtkAHf/NxjcHmQxw47cZz/LOIAa+whb3uak+p55
k7nD5vtqrFbDHKM+X8XSCXqme5H6Dh0cL6vduK3oteC7qzFFYDTofvw82u7dDG1D
h2t5ZoEpxZdZZMPJv1vP7cSPqmBXBFCyk7W9RIJ9cLgVpIVOGl85HXHbWpCyLsOL
JDDGWRxfMTXqMlUNYd4BdcnCJsj3cZEGLGTwfsHWseG0Utx4M7HQrpvKSfhxfkMu
yoFuClWuCD8HZSemD/AdgN2jlVDMGdxfnh3BbEgJEH7rghWhE1P4L8AaASY6OXKz
aDnfgEh5OQtJ89bW6vGax1lhcStUMviGThWpqhHzZj07VV00GHC1hJ/0cWeQ5tPg
CEsVM9hSEHQ7OEy1cBsXI9eaHwbxUtxpnTWKw/gE5lV9zu2PiAOckLAQ8rbbe3CK
YJSY2/3xBnuC8f1CM3xOftKQdhokRiV2OMsxVHyEPv/bJrsQUOX96900ZtkIW2Wc
Tgb4gTIyy1YUNjbyhQJnWZLnEUP7zK7JJh4+i0GuZzR5FSdVyBx67XmiHrhGh+Uw
IuATs+xRnHxrdwhEY6RY4J/ShZSC9MjtTgmHR53Gfg5Uaie7c3QSqoFxPWuWUJuK
nLzEFTX1kgQE73QPHS6+SzoByeA5CEgS9Bs7HpMd8ybfXMjcJCFGOXMZ0M0KPI4d
P47O5BRf82+cZoP2j5uIqV1l3kfwbU1RhROww8hI9NP/tlB4HqVmgR1aPToRTQ+o
+Zo/4Tku1qE3bZ6zPxNETrAkFN2DR09e+Jvmhs7nYO7GDe/JjGrWL1DTG8NbX2HI
swgROkpnnnEN5oPzxBFQLUiuchoANN5Efr0f5wx3wszdqBjV/JS3JCHviCL4iDZi
xcdXqalVT8uoDS6fbSEZf26k7B9RTNr41LGeFUNkFXtEwx0QXVsyYFpQbbGxDxju
uFopnRsFzYiJeglLY51Vrpysn0YYKViU9q699lZZKyr9BH8i4zlcaPg7My5Bn50Z
HFWV/T40ViEBuJtzQrmy2ZNxFolIJJ5SFq4p54gK81I6ypikRgohGlb8YpyCA2g0
Q6Ew1LlkqRbN0NkWfxxbGZl//OkwroSF84oWySvgNzJxt2RwMjLg++zDUevf01ot
ZK7IHEugu2j8ofUao1rkTBR6YUsA2lCvhyVQm0dmm5g7QvsLppHO1m13883qYTUH
LrpG5SxDB3eVA/BUH3/ZVe3eT7a4Sc5SLqizMvfbTqHkY0gLldzMI9epOx3wftGo
/alrJrFy2fu+mEEJA6td9Nox9r3XjVeqRdP1qYsf7BdGk9pJvxDeH2OfI3+R6FRq
Axlr6+68lkFq21BwkahSwZNDw4MwyUEwepMoTcoZDjWvr/SMv+Vq6/BxX3UoxE7u
ISjxoZyN7aUn0YrpSIH90pmi/dhu4uDfZbRub+hko/4J7ADoLVPH/Plll/lOWdu7
w8f8wF1r9H7TaHRCu96yErjAxILUDvfUHTqqVXquqEAIEVsjCLKmJVVWijHombdi
fDA159JpVaa4e5VV2hvEAKqLog4Qe1NBYszOlzTrbyAJWwT8EriyCzZWixqtJCqg
7HFieI7NJ8dI9ppfG2ufW5JOAVV+dhEX2z0v+5Y3x6Wvhy/sn8Z4X3jtawLhmBee
0FtAXNHpUCOjJtTqbBH4r5pIrRSArcDgzNHOveqrgMqvog2sdkc46EhYICvd+yNy
u4zFSrv+LKSFBXWiqZRFQlFegdaeTKjF5frZutZ8vTAWv1Hrd7aa+SntE0uXc6M+
+LF2cgE7I8QVpKHf7gzEAJbj9KaL7wetNljELymjSVQcmtdyuq8uAiYN09yYFkn+
g1JQeewiEG5UciiyjROv8G51xVvC5sFtThUr0td3+AyIAwLvDwPFYsPdgNmEmdt2
+j9LWu1OyqCNlOkCfqiFBnVCIIJ4zWD8wZA+n4GfdthzefwaXOYMlChXiDplezVN
7QBbiAQYvlzltzTOG7nXGK37hhZw5lP7aNYsiavPwzvAVc0JHC7l7ufyZGAoS6OW
jf4nMXuOxjSq7ZNwAUnQ1sGo2YtzzbBuC450Af9+vhmcGYzrYoB9CM7f/J0g2hxe
OTXKMK3tN2ds4lOKREFIQRKyvxS2YS4382p8cg2MyuKfHZBYEmGkYBNGyfehwZfT
68ht7az7VjB4t2Zk8U4AA/lWAR4xZ1ljVVbzkYAJa+nLTuga+UrfjthvrWCMQZYA
jbiMgax3Bc9OqoeOTmJWRmv30LrZ+I5lYQPYge1Px9Snx4mmYFWJZ6zZHJ2anx7Z
UaPfsBmCutjiCJWI/p9IMMJZLx8tfnBPVCVB8UKNcxa5p/kTPyELio5dwQE+P+Pu
KhHMy7rdZr3zhie4Asnd+I0b4ixy2eG152AYW8LiP9qeHkMdQG+Zz2Ug3bwxpZPD
cmwXrrk1E/hQQCqsPtOOnSd3oY0uEEN5u4OC5SIoRu7oxXlM9SfNRL2ioauvIQvj
vYie/ehU5n78Thq3dohiugZQr/atWkQD7aQYaagR514vyQG+QAPfTnZUqZp3EWP6
JScICB7f6LY6GTQAqrLpFnseL8Jt3wiV/0ozUO7BNBklgxJDzL0Nls/u2INmRFIm
YyU0AAs5QEYqAPUEBaEonwApPl1/ldNEJRRHJ+O873ZHQzakvgiW9dWh7sE9V8C2
ANHLA7/NnaiK/v/vCBwblO5RFC8Q+br306LiAwyahNGEWPCDW8/xU073+N6bieXG
L9BvDvhXy8P7If3qr5G3go+kWZV9iC7WCNUZugt1G+ZYQjoaIR0ikAjYHVNwZ4Xv
mh3a/VRib1i6yQAgthrZ72QVIrknLCZpraQFA1ix9PXyarbHwY/CumSCqtoZ2NWB
XaTguA7gWIBEi8sWdTqbIqvefivSz9kH8vecMWMs6k8R5scWWFSRFqCkOQya75Sh
vKP/4M9rTghiWV19YhYpI7t/2wgqNX02/zLH1Qd23jG56C3mSWSvrNCt7ypnrCWJ
d8frGsmmLL1Plx7nvWC90NZ3ROKhCy9MzszZZJTfh7O+KRMcNWKUP8Hp6Eau4UJN
bF1HpjfHt9hHkjevlJwT4qmwFPheAHE1htLQJ/ivtQHn+Kp4PTyeI7ukBBTMGcra
tiisZ9lqT64L3kYWe5UQE8f3IHhCaPD/bDK2zLtUXX/IPJbgT2hBFeLjdvPGIaMP
g5XuHJtrxmiXdxpF/5i8yJFNIyJNiRxFOr+1k77ghiliOhjvmsaCJCmSDsa1BsN/
M5e0N8O6GRMm7fI9WUf3/CtDMjivY4wsi314ont0Zo3wfg+63EEINBVA8HJ6zu4Y
VU+IIzdF5gMtkZQ8z7Ai0gVkkUncOxCPaiHgofSwbBngbKe2owmB8vz9yJUXM87O
KTb6+2OgZA1b4fF+AA8thX7r6Xa6VM7L9h7bGXFCxOk4wW5TC36yQ/u8agQnT0PR
EYSLGu7b3bC6xspjfPYZKeCfWH9VWB7M+0ErJFevQdOOdq9e/wnQm/cTrVytifei
w17GyIOezqvCcWeB2FJ5cYdgIO1LwGpJ3q89etnZImyeqto4djxaP+Oh7Ghni3Yf
0w8Uj0uEXbeu2TuVwhS8EhkPt9QS/UXZUshrwRX1xjKtwfy60VhNPrR8B4QkRAeV
0dq8vU5RcpKbeeBVRW6kxtOvx82hlYlaSb8soQGk4Ld0N0ehskKDNBh46mkXlOzW
fAvD+1jo/mmwcQdb130GOuRLQR1aSS5C3KGyUey4ZokglYj2ErmWZ3JrSBj3dkhE
bSB2OASjVH2jxPO+a0keDBK+1E/wEGa6wwyc10c7cuDZvVii7qauKX1SXxblSikn
lOjbEb3FPB9mvXk5XeRh0BZstaZLqGi+6Pd3/UKpvFS6/1Isa2n7mN5jCY3mShrs
cx/CwzJSruZNk0NasbkfMTjJrs/XXzM9DhPqxKG++e6VmXX5uqZbDAqjbHduIGqr
kGxe9as0mKcvsasdqFflQYNZHk/7O4bVbUVI2R+pb0H9abvKJHun0gTAZJFIXevV
U5RVtp5buDz8h9ouJ4nDP+w5jjtRYyztIbgF3eH70793kNygnzWJnlXrA3jEdl5V
fdUSvYWhH00eZxsEf289Gn0jlnPrwst2LGVadWLf0gEJwQgiqQd7LSJWPajlOtys
YM6uVIrBR0KE2yKAC1uhri6hwTUbpV1Iq7HgJOlQRm4NnPr/fBQgW3BM0ME0Olmi
48b+VucU/CT3A3VQKEKRt42XbXKnKkuUT/RDxNIHaeiWcb5FIC6i97JLn1MDRzf8
JVlsyqygjkENiwBoj8WxqkDgdSF466NPBRBgXM52OtSDYLN2UVf5/YDtY0rhZGu8
dr+v5jz+6stodgOX8HqsW5sOhPSxOVOABWCDsxC43GRQluEeFcXBg4ZAQyHcLYPp
RzDt3JWejgqKHi5OShbleEeLbr2GTxKxzJ5V4Mv0AgiMNVSDmEIVdtASb77osdf3
LwcWMW1afDUkYWcg1hj1NF/65Bx3PaC0++xHhgfjPGBn2USh2j60ddrHJtqqlzBf
M/CdlWcFvB7AqD2x3lDrKwAWLH6JK5UBxUSb8j/RGxKaYdyV3TTL04Qh+7mluKtm
uS7McwEfeA9enFJVlunQ3a1y/JyOCoOZUuHH9sFQToze5GCUNGtH/jzhhbRIlydC
purNJ1g5SHsubrOZiRlYOIsigHCu8xB1v+nEUsT+2sc8+lazbBBFMvlXZIT7cOVO
oyzrJ+Lyd35JoL09nk7r3+88mlgAMn5JuElplCWWyFvvoQKEM7Z02qMRSug3q9a3
F7g7dFmW9kkto6uQyWRpsBnk/jwjE4MzEXyVL3ZihxI+BkokffYfk3af2Gvbo6ec
R/Heec3E4TrZl7IS0SNDWKdyPxTbmAsaibnUvZIk3/YxNHAqeNNwLy8zk8/32Y/s
OK5tPZEhMeQqUDgX+sZW2QNF9wQydrZHHgeZoZm219jCFO5DZ0waKJIVCfxBobIq
R+87TOWrlBBnhK2rRPTjxLSDKZsOhe9tvBPlg/ipVWhV62AkzH0qhGCA2iUPVU0O
bqntsg4L+ZQMEm1NcsaAKTfjRS719EqGQiLEc+lKPFSZKrk/iOdS1Qmb5K01VWqR
Qr34L1wF8CLhF619Lup/r+bT/Gyv098TerydR5OV7wJ0qVItW+55va2Q+zjokEjb
QxR0Jwe2nKUY1qk5VvUgMrz7lY3iU0v9wR6MwKZu9vPr+4Ixh+IkFvRIVCD+59P1
gU5lWcSRbdudxhrUfbeVzdSJahmKAZwBX7aYUb05u8wDTUWeVL61/1taiqad5x7N
kySKIh9QKAVs2E8ji36wRqL7Ng9xfd62hwk+wwopD5tBsL91FkE4RBiFEQhBlpEb
iIZ71Hj6sl7HCxQA5M5YFhQJJvUlQ+5zLPtleAR4KBGv+Nev/8SZOTQQXI3RjOMh
/1EHrAVNgcmLmwxgwPJ/E0V+NjgUIQGw7ho00yq1z8memMctVXIX46TqMrxmX5mD
7souW5kHt2ULtwEbxqsQVKH6d8FCIGxC8c6JWUx0LKzY0p7dyMiC/pqMDryiIh8P
93NZyv1b+nqDaXFV6n8xIFeOfOuXCqaBgxRodGrB3ifD+I4bpNxiyidMx66N3Eud
xjFeZl1wCikKb5DyoOV5taJ/RdcbFajeTjKpEuoMcKmaVtQY2yMgpO3L/NlxEt5V
xTkh92hwh9r0VlR4kYJ5ZQiAOaQFdONxdhYzXBGoRA0ArIzSZBw7NsnYAUTFRCCJ
drMILjcnuKrzs3mzvdg4jKXDuqIc9GQz3U/rA7peYtlZ9UONW3FWmVymn/SILpC5
BAtWQZvK/UBVI52RGEh8u98gPPvv3GP2+0pmIZ1nyEvmw3oZK3x+P7wnCjBDMAGq
O04PSfhKlGYfkSzfQnh7zmQUKLHVhLCcGyUmuzfCPMto+Q9jPhgwbBf4vFBY/ugN
+J1Q1Y54ZIoNsz5xVJW3scsVbwfrDk5SglT7Oe0wCiRKGzCswSSAB+VmnYdz/imV
a+JLKa5V3kJrh3MoWVugFTjTbRgPfbxHiLHDjxbYdPhziWoZqMWHa2ardbG3Z/gO
+NzKsP94dYf93Vir4jtrns8bEyaNZcS1bAh3fUrwy22B4CSb6jhLZVVBBgxShl54
3aT7YJrvgS5ew196TEN8fEaXezpi3YXI/GHj/ZQB0nZMObO4R7xUsgB+u/eemg4y
O4vuiLbPFn6uO4aBG+BFHRqsIAWZMcVKb0Bqe2GcQsnCGXRlLZFvyIHQNwtMRWaT
U6Mmpa2XAv3vd13arDP77zYKixpZFpG6U427rE0m3OSYOgQjoAvWbw0n89M1YxaB
rXFeUT73k9Uu5UDcBycCQKvYKSZgsPxWnvHy42F2z4O+dWsbsVt4QRdTf0gZBti3
TRvDUGOUPwaEj9tw87obF1gmXheGPgDXm48urB/sAT53sv5Tiz+/mHbGswQ5096e
LPC75Uc/QwTH90rtwYj0BI5fWtHwOzjmSDQncsJ4+2T3REx5CnB6QwqNN7IyQ2b4
Bc0cvmNkX9//acmULWQWPEZt02K+iIp/qDYFiKV5ZQ2uBD/DTOmORyGG/hkttVXl
AMgUPAk1rp8pJFOychpvZK5pCkRtf0xLfX+udsPS1RfQS8yvjB17e/7rpBwoohoF
biRMwI6gZn1zdM0lZqvnAXia9jzI469aPZZKYQsC6e6ZftOObQ3uWiA25z8VzeLP
DBtmu9AzfI4VN2NYH+wpJXc0MUiLY4UjsCzUtx1WvrvR5YF8/FpsDMMdF1HBMz+q
/cbBCPXzOCp5Mq4+RYnMGNBD3XDYut4MfLRThJdL65lNPyCe0SPqrycTY17Lf84w
9AH2NX+51CV0S8lM3oQG1ZQVrlcBidK4ATh7n78YM4BlOscM7mr8rLQSVs2xWI7E
3cdl9GHrKVUFSnjxwud11WMOjAYF7kXGhJ60ZNYCVcxdXquI9z9LRkWqPcIRY19e
vj7s7ov8y5gjS/LPnDDNEaWAzKBgw9/mvcZC/0+k870oO0fpqAJTvlI8yoZPmMvJ
tWyDt0eBVchAuUAQOHVUbC2NUvBZPr4jOiYkcrbDw2/grZ05rBnOH+YKIP100haW
xrLrwBqbY8ZVWFThqv8/gAoElPSmNabC4NcgixlH9jcmBLyuoN7tvH029QVez4fo
YDKisIjkqh+OBzrEKSY2lZxVY2rzPTk/Q3DrwK4i9hCeUgNS297zyWyUCb+hZJCJ
LQLSrcp0SvG6lZC/6hMM0xc+L+hg+ntegXOX4LQ58s2AcwKfIKwvvlNFLfhIyIW1
DnqCleU1oxodxMDGzBHI2RADC0tInLW4Vo4aSDtpX59nwlCRVeuxsd/4uJpfyfSp
J/N1OV12VS4N95Q4eFDJy/7xfURiexNm/vckS5exd5bddvXdalRh4kv5miu9tgZC
`pragma protect end_protected
