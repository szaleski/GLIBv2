// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:44 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
AlSSFLijnL9CP2Jdg7O36jXHleMGbmjnDZGqPqnoqFBtp6M/bg1Lnri04d43/1Ep
zWB0QTjkSs48jPM94MqfSv1EX2N1SI32OTjegmR9rpW/+qybJQsjAePPLpU527mI
lljNU9ekKGg8WwxVGSC3QXIh4sDQoKyUjJJ1++Gh6SA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5968)
Y4e6UQ79bzvEY1L8WgmF5VK5nmGptt6NbXt59T6OCT0mAZIPre6Ra8HjdHlArwdw
ECmBTV9B6+/2Seysa1vXcttIyI+zJEtKTStCfACk26wGeN1DtINSJWWSuavGOBSx
svVClvCYCs8EELermo3UIxWep3Ls+BCY0smIzpcxk8o0XO0bpggKIvLlirS3snDV
HYR6UousqTR+7Ob0uWIWnDzI1FrL+sV6Pd9RAJRujYh+YWi4uOfloATrBJV2HOoi
nJ+LQPD2S9ycY7RSkUph53YjBGqCUecl8ai3ScqDfUiyHV/5oLyfx7LfN5aPLNJZ
kXDCKwYylenePpTLsoDKL3NMXO8j/WE7y3q4L7YlgDZqcA4DtQNnwGtqYm+D0vFa
x764/wA5drelhC55maf1kKiFAYcayQde3E7oqFwEsnNhO/2efkapK/YfJRcSgAxI
k4ZSffhEdNrOhqvGUWq8YgVYoGVyzeiN7Gr8xElmcQ3dsrJrIUEVXPgMDjUMuWl+
q2JH+czstfL4lltiBtOD4b+n2lply9iDjKtmBKvI1cgqk6/mkCw894rOJeG0QMfN
Oiwa0RbCuRGWQNUKH6CgK5pIMF7I31Ef9IuAFHOM8r1zAwzfezGTRdlQUyQVRe1w
kapI5d+WvOWQB+nc9Jqout6hT54/4CSUciUU+TKRwFNlPG5Bu+wP2ZYpnl3RP7SI
BlZT1u8BwyIbB7Ps9iM4r6vtdKtgqmcnhOaK3/AhkAm+YLajUkGYNEqgbGoU9Ltu
BbekbZvDukQWsgU3xa1XZxFG6QduIQNC5Qb1sduzrs2xXccI0ziEyTm9yls+k21y
cMaf67DUZNaEwGefhEsTN7k9M8tYknPOD5acguBAi9+mTAwsH/v0zdjQd74F1kf0
63rUegfhgqSYA6fr76srIGS9YUKLmjT/lOo3nlu4sKUjO8rQ5fXjz/IxsF4zoCF9
9fgi2HBPkgwVeGCHuDub7GlCNDBblVVpAyO16gQSyKWPK5yeHDxMtDUu47u3RSJe
S5omx+EA0uqyuV1bdWWz4puj58XqgPf8JhWUBf9+jDoxT0UuI7vfNEh0UD01knGj
5pWv9nviZSJ2UqzhoEGLxa9+VTx+BB1LrwU4TWfyn9n+4SMZigSF6ZssiP/raUBa
//wWeDbaWImEb6G+bEBcqcP0X247sMnd4g7whMw8BA7YSrm+raZjd8BRifMRfqyE
7FCJztPvvR8VSzkHVntPnrVt1nCk99trVly7F7h6wnWnTCEAHDLpwCYBRHubdyWV
X4wj8EuKwDPFg56/b4ENsWmEuIx62l6m4zOn2PNWIWxU0Di80qh5so1cxNqB7opj
fbG2l8S+iwgrLZql31hSjRvZbz2affYdZGjBqg7TrpMF7Nxsi1U++LxvCUVlLFLd
6Ru9joddCM0AB7VQ7k30vCcSkpfqugSmq7JqukX8S/TkYRFAbF+Do6auYjFCVft9
LTpTlRirpfWTsfyi2/500bNJyN/G6M06o8KHjxTej/B5JgA7ZYY2jIHhn+o36Puc
GS+HI8VmsGeGb+oG3qCw1jtLi4wY6Dku2DD4LzMdyKCZkPOSsDUxyuwPIkEBbowy
ucJX0OadNIupmisBbSKcnypesWLi3pbOD4JdV11YaP28XSAwzi6u13y68rDEj4d/
7UCwYC7sD/kaxiwdhDT8JlXBgwDi9Gdj3FO6BYgOcVj/XYxjo7ong1GX81YdEeiC
/9cnJrM/sVS4iv5284CzBZFKKb12efywlwEhcEiIRcLBVPcGZaDvmSUtrLWg41j6
FcgxLq08nYB/lseK8XgGp3XDaJcCRrQYV1CODjny//nuaWRXiI8XmTbH+NbBnqDW
wbst35NfXXDlVk8gm8dfluVE7Jyu3Q/Mavrv+giY8zz/pATKJW+Jfmu2pUoG5bMp
2JAN9GOGv32mPQWmpE+M32p4jSmA3z+jGX+rIKfyviju1R4Ej/rAs6Z/L76Uis0j
QVbtuX9awNgD/ilW/L8JZWh05wBlRRuxWz2sH+Nwx64ZN6/em4HTj85v9HBsiVgE
vN+KdyEXB6FdnIwjs08yaY/yjNFPdOEMQoZ70suy1hxp5FNTHLLG5NEerN4uQbVz
s69ebsgli0yILNiOCFWXhzr9yG3mYuuhUpCzQHm6GN5lxwrT6P/3RbXy7NOdlRQe
/lD0qmAwBeuKQiyfgcQpR3s4R6xfOle5o9baXHID6qHJxCr5uMB9/p43D/oe2OcS
t4B1JiTELN6SgqG0qeeVF9O2I3aBUj8BDBtrteccqHEsSh5WBzgO43oeY1tYc7xc
3P5ACCVkKw9t7NjyDoAlqDn50aOzsEJt9V+ZdWNpSxb3TtQhQT+93VNvFmLz34Ax
0ZCS8qP1BBT06lD8Ln+rH1MGKr0FfSFFJ40eTUlxbQEU9iZEmPij4bzu2JWtaQ8I
sp+CKOSo+rtLcu8K13rASWwfK/mH44TrPOirFkXHll2KnPZNYH8sDQbLld9erRwd
wDrbz8utbu9412WGr678lPF+rZe5AOWykblQVTN69nRaEyZF7ZpEtaqDe5/r/zSL
ZIwohpLeu9xn3PnUEgyR8ZblY/zuHwyc032/QzMYM38VqAvyQltNU8DaZohP44sL
83rspD+GjqM21+kDVifnBNLQqw22u2Ac/VLZ7bv94einbOQuMsrKguWlrp/tJF0u
smO1t+aNeAbpnVJ0pqrlT1z2YHqBTMiZSUtgf8BkKpTryCaR3NE6hsmhV7TCrm9W
qPGvC+E89KAHyKWKT+duK0eq5vbKcGqxFveFcQYs/1MsCPYAYLQAoV5x2yBmesJ6
hVXbL/Oj+TO7/iCMSyOex/T4cAGAV+4RnbEM42KTt6xHW7QUqFgUojJkjqn34CBN
uxYsmJhoxMJW6AIBn4FZPiog6fLT9D6m4WvdVssPI6FwjhAhxg8mttk7DvDGGOPf
X2g5CbfiX486NrOquKjwRA/DOzhHfWxdKxCBuBRSTXoZmcDYcy5rRO0fMxjgTZ6l
wQTMEYxedEKyjPV1PA7y11NAK7M5vpGu9jQBkTj6j2sB3DDrWvcdhyehMzGcsn4g
Xa8yDYGMpNVtPNmrceXUtkL7UUNHyNPppswoL1Q2xYm234ift4EAzKOZVtwA27yL
MxdteAgH/k1/YTMRJdE3QMns+CFXbuJrMGgSYYzfrJ/mZy30ml7G7a1Net5EAJsj
genkBTQ0NG5O9LhazD/qZOvHsZFSbF9SeCVX+7wpCK1jJ1ZIhbNV5766eWhpER1J
ahEBkN1iyxQYgb3HLO/xBf0daaDPvvdBByemWAA+rhvOav0YfkbBuxjKTKv88x4k
DIy0uvYzy3bjqLVkH+rIZOuoJWNdYP2ZbRUOn+ft995SxCbbPrrFkwOpe8Er1bAi
+x/A/q0t0OWkmmpM/Lwo5XUobUf14NBjobjej4NbHCXhWSgV+Tc0UyjMRQ+z2O+e
ivzUQbiW6GAV/2KxSEPF9YpfHaOtAo5rzMg9c+QrXM2UREqWTFCItABlB40+pZnZ
9Fh1E5lBqINP0lo2DVpWpG3g7oqvIu9YCmSz+MfadhFUywlD8+qEyk7Sxkj33++D
wOIO2Z+1DASaTKmQmBheEyzkaCl1WNzI59XJIoVmoyNwJ8MsfNzMP4Xj8YxN0cKm
TLNW09j8UkamKCT7z0izSO54gxHFlVsnKx4s8k/hQh82WutbHx4jRtOCebf2q8+u
E1Nd1Pg/CdO+1s+ahYRhrZsY4l3xgEB1D6/A3Wg3ocTaDDpewvateAvNqg8da9gZ
UX6aUKmc1GjKAXZyKzy1lqJErmm21/gFHChrnDsPKc9ptstwMsz0PVbCBK39ewsA
Esc6zNapkC79SdJP84c5eihpLEqqYD6NHPqw1Dwl73KjlKbdeWtMkplDKk7MfsFE
DZnVj/cY7Aif7dGUzB9HAevwIPeOQ067nNUr+zQm4RLnAQkYVF2PGG6sILbluRr7
5WuhS3y+XDz24TGg0s49Rpusig/TlkXWhDEItc41R7RVc5oO3E5gIkAXDQkDWEZH
pLmDjL5h6sy959yCkb93BN+068w76ODY8Qq2laob4ImQD4GKVR+KSmHHfBDBBEq6
rAIUqrx1w5fzhMyxAd76NqencYR9ka5IlJPH0ZEAlmN9LWkB0Ht1w65CYNbOqDpH
SUUWsOLKWECn9Rou+bbMMUL0A81Tl/9FkTrdHrkIwz8o5yDNi4ErjxkEglNm/67o
9mnRQXjd1wpH/22Xg+RH4GajFymUzNsvRF7gyXPwZuruMk1rRLZd9END4Q+zhyBf
ZZkXqQfUIAELQ2Alafp0YloXl9sBXkAT52VN6Aq0zyq50oBcm7ADrDwAU12jSPpW
qQOdy+kPwORGrLTkZMJX84A4KXkNO8ZsXFc5PTtAtXA6nzhSc64jEpvfaK6vp7Pq
asqujhn04+c5/ILbNvrOHAG5kAzjgjBH/x5jbruHK+23Lo6f4viN2MGSXdRsL0so
JB035coB7qFzOgE7sC6OmnQbS5h65jf1LJELFqOt1VqwYPt4aCIxq2oWyontXuRy
PxKXc6XtxkBU8TTF7DlDmkc/HwavF2dS6kCaIOXxCknqn/zQy9I9/59pjUJrwywp
MA/Y9AiDi5wJ2ASBhMMAu7/yQdG/KTdaZOkdbtVlocjEFKmih1FSQeiKpVT1Se4B
+4df6d0qRQr0WyxZ7PK2jZPG7stQJLE7j8+xh/VFvpVUhQpAH737VPtetvkRd5wv
odyvobeqKs+8Fx4+TQ0hxdRFyqr9MkdYpUE/u6QUovJqqUZA+ThGNFMeug7HwoWY
pPWeK+7qbECZmBlzSuyZUuIOhT+Vyf2FXW54YZ6QY6m+QkfNB6zrBMzgv6Apy6ux
m9tr5cGCEtPmmBGyNSQlmFiMhOLaW8/I9mMMAFDl8oagQkxE5mOgrzLjkqma4APJ
JkvO6Nv6ii6MNgclv1qk74QfCIryptIktTJCyMaG80zFEVbEp65waRqiI2ufKjZd
P3FbC9vm9SWjTqk9Opgb8SjKnkjQrdWlaFo/pyo/Hbo6mnIskv+QJPHi53Enft/C
a5nM871PZ3/xF0bbB84BEv4UsXdzpsnYfx+LGQdwbS2IIPZokKqJ2DiqpLFQ1aOd
X5qjVWbifIl1jQpY5/a7xt0Wg3VhMUwMKMsDHQFZM8V1LOj5TXZXZU/eC66hsHKP
KaefWh9Hf2uaZX5S6vjM7VRHuR2cknELptLyTqM5IWKzpo6/sSQEPPj6X3jbILxo
lQjLydFHKRgdlf/yMfbEqHGK7lm8q1lsZsGeJjGtPN1+Jwjum/KkcNwGtbf0Ig3U
kCFYF4G76oPqCtNIxeGP8EpLk+AnpxMQF4F9hgR1oDRY0KOh/GZt7CjUvK3uTctn
vDBL3Yvr8sRfD8WABEHIxfgir7ZzY86WHW58CEj3N+DZehQksdiEM7Kg2c1HAr0g
dvkS80IKFE7knw5cSiZYl4XW9MBwVIUVMsPFObsjKm+qSj73ldKt25zzD5QoJpNY
KuByLpDIT40XgtZ6uEL0frJ1F5YMFq36hhg3Et5QBGAnqZQdvMz4bgIJ3JEsQOjk
muYYIfbVuVTvunn5Twr05Tcvx7Axez6nuPCtpSI9+4z1gRB6liu10nWkf8MsxiID
cEahYIh74mVUS/seMcRQdkCTtmeR98BGVRgxp8gnBTX6X8QPkeCRa/JONEPv/I+k
JBnp8PsZH/lbgmLJnG8D55vIxmyqdwzsM4TRftGPfmwbYQbr02wCKZ5jhRKLfzHT
/3Ad/parIaSn7GguyAEScugzQOtnyYRF4xlMnhb3Mx7tSt0QH7gES7reja428zCB
WvR61JDnGUAVAsz1Kiz+Z2yTpjWlRW8og81vhUPBqscVMJ8XcJ2I5cNclePtDmNS
hZ+Vz5v3e/jhNMeLkU+Kif5KYMRlVd0RL1rBEQzgOvBR7i92ElVijIJIfELcKOt+
M1oEMM1ZNHsI4k6qjtIPTI5EZMdzFyERTe/mZGmdsr0XBrb17RneAPVvPCqNoEbG
R87LUfNekJN+Qd4kJP5jeOdnQ6XOcM3OC6CUgbInoX/TjLFeG2VM5VHzXc+mNkyl
frnVPtvFufy0Ya2IXauCRqrJ4KrjEQ8U/gPWlX2WESgskZaIAhn4NIzIGX6G9G9g
ub06Xla9n8U0RfL3LTkuPtv7OkaDHCicMMZhqWIttVEcp8biwlt8nO6VP2Hu1G8D
GXJAQKwLbdf79EbAaWt2Y0BEOqgmMOBGboOx5LGTd4vQiPHYGopHfcB2CREJsuSy
zIeSCvA/YVgfMZKPw0BKFFdVHb7TityqR2gf6yJ3mXx5HQDNeEanU7X+joi0VcGu
bKU2NxZK6EUmrRNaAoqvKqLMq/phs5vscRx7LK7NtMYgVGldKg6K1LnlEWdmZcTL
LxV+zVsBFnFnfMTchQTyqqmLuQwMRWtkHBnnjOap7G/kqjiKb6n/Aq2gX7XhMFaM
DTMF4vwVi/GyzGGOMRfCtDcrIYrhyoriosdb9RqvI/MHL/rHLwSsNveB6ua9IgpO
2ihNK6SqN+CzhDWOJb4LrElYKK3YzFTNYJDE7uO8V3MnB3IrS7IBUKGuAa+JGY7j
SZ/N+mvdrmVNcw5in1r9ucDFD7k02vNnPzJit0Qlt+R2fe7ySR2kiNBf1nK/PLom
sK3oV7p+IEovcgmNUh0sUgpikbDojjxq7ah1rglHpXtO0cFYYTY0jbPi1Vhd/8RK
ayQ/Uk5EhQTAn+5S+4+A78+dOa0bcRTTu8yZgjSbUbIP9ohHw0kVhrWflkBBvqbc
QQJ37E/Hcrl3+AF6XulMEpMlxSBz94JeLevILG4Q1g/dDCx57K2sjCIAazSsxN7x
83GkEjkyZK0LK0Pw0wMqIpFucXWeZLXt0Bfjyy3XWUivy9/AnKPr11SFPdAEWOXq
ut0x/RJ+0QON1wkBLNTw2rL7+tgmcytYLD2ihemNEBw2EJMJxzIW8wJTNJPtC1V1
PVj7OjQzQ7at2+x8twtZPW+nV1UgcirjOICHt/PdYvpyJG5xGinn6pCQoiBsUa7c
1C/DWF6+5ST9s5fol9PLQOe/cpJEq6v3YoBg7RkNODUoJ2Pb6w6r5RbHP9RBZopb
/tdIAohECeqvnasYWHxZ0/FMRS6oDDBpinJyTSYP7Xfa4V7brrgCpbWpBwWWjZY8
o8phgrzi1KMfNgk14ZTdIgll/BCmhsYE30DqKm9K+kY+osCjYlqF7eoJzgWtkovB
bCQtPtP1U3+qpCzn4QAGx54MEtPB0C7gTiv/BeJfFrZqnvWOAfHTdmsZ9+DTQKM7
dGqsXloOjLnvF9BK0CeBBSx8LEjjkjoBA2uvzEkoClEnu8b4NG1q7BusZwF60dfD
tscNa7JXK70H+nXWxGQ6Kh7QjcT8FF3oohO+f6lDzNEM+0WDUjjFA43V6RHGVOnx
szeAC9kodlbi4u26ZpstiswDH5hliGHaQaFWfnw68MNdjDJ5LujKrI6jBvhFg7fv
DxhctHu8HAC8pKHghpW/8v3evpAU2ntAzisNrXyIsLRK/HS3OQ9aon2ARIBE+cpa
4c7Vm6FKeP5vpUhxMqw5J9EfWEjzsPeiyQNIXOxriUzzZ8LUekbFdpjhjOyqTjvW
E/XRfKoKj+w3a+VNW4A1dT3zy2usvMfbyulq1D+3in43F5mRiaKxD+X76wOxmOzW
U6ghBWryV/CNuAV4QL/gfQQ68CNrTmdjKmRfIBLO7ZhHSDYlPYttOXrZn+3eBeyc
+tr0GBc+rf/vaPFlgv1jdj3nNJQeK8Ki0m5x9TDhiZgxfRyw/3mTNf8F5/bJz0gH
2tCP4bMB+ZLH1go9oxdj1kGQfj9HyOIUqGPyeebLJmQLKxZpVZoaLMOWubWysVk6
FCeDYGoBLhJ++zbfAMf3HSsR45ZcWw6poqB6gi1r01wjGUoYLyHXdfScqu4/3Iq/
d39lDMZw5+IEWSI1Ezt1SA==
`pragma protect end_protected
