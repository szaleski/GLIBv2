// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:33:05 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
eXjFW0HmNWLC32tnTQMFrCLJx7t/xU0T7r2xQ3G65jPWmnGrWkKsuFrAB/LHLt4P
uzbAIA27PnKmT/JSQw5v8aVI12HigElco7U+wqcsUbHySqD9Ehpo4S8YfgivZu9T
ibly94y3vgh09RwM1PC41cyZs7fabwdBshh2AxHeb2c=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5712)
M4iTq54n9WkKB+yCzhEGOmAKiII6hWzBfGLg7wdFBBpevmi3o2Yvure5WLRaFXFj
LZHuUuatQhrrLOH4plqSUQQ8LvDaBP1nG+HjckOJYNn+NZCw1qNCkkm5Gkaeaw/F
w/4iTGnxV3NCBKi7sUg/SRkCihGZPaFaSZDcC6notGh9i2/WY/dxGt6DhmwUVmul
dRh7qExTFDIjVCvjkfijxs4l3XQVjC8A5xx7x3tWFmAmxlTQRlxNdJArY5VDo6x8
js9WIK/ii61W68jokNDLcHPzxctvK62lAZ/nGb7Lz5PLM1wkml8QgX7+RoHKnc+R
FszpVLjtElgc4f4Z2E34Ca+BIxPh/jy2TAg/QZJaDqiaQ2TsuBqPTSu+uZX+RQhw
KfUX9H4nBDkjs5mI7l0bVNOJB5GHLXU4p62KeXZ5ew7cdJqyLuxwvJoPB8BLPSh/
CoV0C5NVq/Et7kxtvblaF5z0tbMweRumPyhtoP3OJeb4zHOfu9JpdlZK787GNnYl
1pPWMX+WnO256yNxbRBz8vpUxWoFkA53sJs/jQdCdJZwB7jXyjjjfvZMpPonltzy
N2JPS1rHbh6igyxgO/Eah/6gxtgM/kjFxgWMQ39aVMTjNgSFM3GsEAeG4xEAveMZ
PttMPEz6EeQ3lKmft2oAF7ba+w7L9A3Ba5gG4vNxj2KRKGsO9Qzesy7lwjdHDEUt
bQo5jRUvRPOMSOYjlRa9W0pCqfxpG5AE4ZTkZH7lpEFhI2lGFNJMeHrPnX2CQrQl
lPh6TMjoKixj31+UgGKoOxa3Ftu/KAI8tnwLfDMQtUHUMExuCjHkr9r8M/Ca+izg
yYQMBxyFCaY527l1/ga8InIWoun0Z8+HQUhS1RmNW8ToAr/BznS1jFfr8ZTG33Ky
G+POlLiRZiNKpLFUNSlRG2aTM1+tzcnBKumHq5iE8kvLPfaTHJc+VvcrNztvObuV
iRrjyzLZKfiWcwWhaijEg59uh9FTvLdwZABxSUOaJl1+sINOcVV0OVBOO4pywqFq
XS/0ix8snT50jAWUjVkZa7u3p5F/SeFLSRSbjIXejvWIThXIezFut5BYaR8un4nz
qt9vgi2WsmroL5Gnb2D8fEdNQyTSnzhZTusZPJGhOkLxkxTAOJlCMvuBJUagumEU
M+mHEI4f3YdAn9L12h9VYRWN5sUwT29gSAxI91XmvrK4/cNKZ6JNK+b+RtgsJ0rL
Svo/jHKslAXpQfA8UpPadGke0Uob386rbHADDGJuzwMeJfEwqMue1J9r6xO+++hH
c/ITr7ZxJYoIGD+YJoqbJLmB7ekWTmm10djW2n7EFjQv2r15YOB65X7Qs5QdwP82
EyOxJshuTj/TXqyVuzaAwUzqrmHo1NWFj4U2wOtlnXmvJKhmretauJIVGa4x9QPk
XPIbgtaoa+B+KzDKHdhqzPsbB+q5LCAcY+3WR4b7vUj4+P81NSVqeLErW8zcMKCp
GEQlGIWv8mTCe9EC8OaVGT5ItyQqlou+2Ls6e0Xxw3EOH7gJov9Sb7acDGcZ3jml
yJzjXA4CFhOH98DQRbz6K8selmgrSf1FKnrLu5HHjUBE+v3RO3DTWp4IyRXJV3Pr
aXxyzAF9igklsnCGTVwLGZ7bTWz/C0G3zxbnZAuyenLZiVfpoG1unLss+3c/kqMI
JK62FtU+jCm2hAGXXlq5qX1XRagurcjQDJj0dwGoQrNWcEVxxxtkhcCW4EFVCVf7
bc8IkwBrM4GPZ2AC0/gFa4qWTP9+kYdibSiHnTM6prVxFRjNuYlFCTfaWo+fJYXY
8RKPLCGeERHZz+GZhksxhX17zhr+1Cgx9mVGlcOouwK+v88COD8bRFvBs15TKIUE
uWZr5suXJjQ1jveEwkwGleJYeZLt/dwBrZWVS9iJhypRZcvOnhpHQWKQjYG+ckmt
0dB8l0EKleQHLNvlQa4gGT/JraH8m0ewcEMx4z1ut+o6b1/l9uDuFrEs3DMoukW0
8QH225X2Fg6s0y5Rdd/Izt5XIGUEBpDRkDNJDaUhIpu2TkxwMR1VMh96ZUU2Bpjp
BNLVV5lkvUw3xRyEvHD4gkw6ctYxFkRrckGlpaxcSU830GneNq6Pa+p9Zpr5YrMi
LjmYvqMTPZiNuzdmq+WPnq6gUDHc/MBgy5stVsrRgg2G2B7p6Wa4uYy9dG9CXMnT
5EO5wXr33GZaBP3Ks2H3Ry+AooifY6+VoOoya+2lsdmft489cnzJyGA0LZ5y92oF
C44QJ4WXcWkNvu8lAW6FztfApm2TGxfP46mLLwTJgLuGscDgw7K5lxOfkP28IO5o
V+4qG5MTXZazgkRX0K/os/oLdMBjtsy1e+X7SHg2NZCqVpqTFkCKSgt8B1ICrK6d
cMulQteKT72UeHjUgSClRB0v8puimTM92M8pIwk7PzZ92LArGkj3o250sh0GSvMC
uzDAhnX9SEYQq7VOjS6v17oyoA+ew+n8FTiYXs93rYuyfvvq1Pq1p58EQ3jNTvdz
bnZ2aO1+v6R3yPcpEVhCbnJZO7OOzaoyEN0HMFW6u8ls1IdP4yjn/1zhKlrgQ0cF
jsXKCtOuq5D0qXXtOAnGRxjeQjFmarhAU9MVUTuhby55R5XVuyrABAukHeaVHnhu
0b0d5a5VauOPFHCMWCT+HgZ7w5vbvLpz+P26/+kp29YjzBKR1pyhodowdRIq/I4W
spmFcdVEdvdedc/N5BmBFP1pfpg2BWQNsRCAzAiFFvgdwnzCWZ2wQxj1kcatXLFm
XcL/kflnF1GaXA+4lXwQRk9iMULSz9MElkkGSsLhtqSOLMx47iGh+ECe3ecE7DeY
N7TM5b+GgX13FlGwLa4Kya9nXmnKOJom+lsYR7c31DXAIV5TCmiL9i7JOyEUJMcO
vQjcyCaNtnPR+xPMWf9hNM31mmJaDvaQhmI5ANXJDMBQWpFg0rA80jYq+pkpuEEy
ZLQ4AveGPRidMjd5UTpRNnxF1WdIGDXOu39WN7P8TLd55KO+DvEi1tPfEPIdAqAF
3+35xhws0GoSXoHeyBD7qQ+GKtrN3Ged++gUs7bcgEL7wlqAx7DE8OTzPROrQn58
NeSI//NtIrGx4dnOTMnFBy/HRPuFkigJ6VTfNO6a77gfjU6JJ/PjpXTmjjlPSfcV
5/pE4GTn9cfFTNJIsCukHGp9QRGlUl5jC9HdEmeT7gE9pcMsGkS4J0FkVWpWnEgD
jjYY54rdIibz5fJmG76IfDmysAP7LU4hBIj8LFK46BQcxPLFGQ86bozowHMRRUkB
QSpJvammq3WSw2glDX5f/NVLmr0HftqQ+mgMcXyd95yg0k3IsTgrIoxYaLZT38C6
E7brsWq3nWu+B8b6WfLFe/sxGnuwJ0Zg8OG5rVp6cKGlymvGAX+lttNd0XoBmB6n
us+2Jp2ii3fg3FxQWfcV/mju6jmyONr8NGqxQGVbahJbsRbxcBxkVa7o2odLslIw
rG4mk1tS6qU8pa8cvibU0ZVBzD50oJjGk1yZfFik49uFDEolxwL4JDKW+NrCz5J1
zjLcvYxWgfwYFiKDSXc2LTpZavS+vL5IGvk+oM9ByVLapmfGcF73Br5mK4NzskTv
DIWsWsC3yuDavaWUb8XHFPKgPVr3E9MEM6pXR/upS6qcNLkWWACCAuT3tt2wncZh
CW9VutKLnUVhXA2AyVKMoAF42HtSmvEy2EfrpEejOhDlD/Sg+ENd0CcYtozFVipD
V2Z7tOlGwAyJ04kRzuOXZkIoshQCMLsUkk7qpzT8LFdoAh+5u5bbVRq4sC923sFV
CDzRBzz3gzxsZM8ALSq152Djt4RI9ud05XJiAsJvT+NtcKWhNu4dCu0vUGJsEXx5
o9iUcbRGvLwtbXrqiCSiWnPoUEf2xObBYQ9MxwvWNT29DnSq7MUFnWAJmh1BPFUX
p/hcYkar40L4aY+pGE5RBCAkY20bYpLP7yBf6m2JOqf5QiMNXg404FDy1L4oF7SE
7O7TIHz6yj5AKRNZB7ivRIA0RDivd7HCbFW7deq07ClaYKBR/J9EI/9iuKjOoHhC
jOvTWJ1SAVS0HCZvu+TcaInTF9eG0+2cqEdzHGcvDdjgpiXkHl7sp1GM7146sdFu
r0Juxu+x8kCZFAnQ9+7pbcWJX4QYL3Z8tFvw0XTUGA07k0Vq2i20pPLkbc9lP9a4
Tu3z2WoQmNsvGwELMhfXhsQjKza21i4oje0H2TONWs6SjdqeOIxXirzU9DSonioG
J2yK5ehQ0N8wm2qZePPQ4SnEOBmtwtpDtjWae+2b0wk+Kqzw4o46jRvFLCIxpKe3
xYF9k86JZLGYGu67eVy+kB0ACfq5MvvwbK2pAEDyhuEA69v+h95KJsjqSz5CJ39x
EIg8L23zr4WyqrAAf3VlgpNDwoaLY6H5RcPwofAKdV1Py4OLexQmmkfZlKu5nGVZ
xTCAwm9r17OkfsDueiewNx0J5TrVwEHs+rclizbNMVr4mqnsZovvdMRukeTn9Q29
vRJl47dsG0qZM4v1Fc63fOAho9xmV7zQbKSGQblE2uYBX8zEsKje1TcwjKqWUCct
qohm1ED1AOJ82QPwMetYO2M4ZgRHspn0rVEY5yWk7K4JbWF+WKDSGNGucwjGZgWZ
s8dl8/pEBD3mJ4FwhZDc3Q7NXNOYh5ytFRiZk+y4CVcT/RaXnNvM5Wj2xENuFMjc
Tu6BgFfRClwi39G6jGJSJqH0CYG4HGM59wlhXQl3qxaWdmaWmpKOgqPDaT1Beyac
/eDUaSux8JvhJBxTKE5YiA7jgLA/wN3nPwGKWijoFM81oim2K/PZeBJ/gttnZbA0
fGY8E0p6lOQY9UJkUuYSfSPWixesmLbOdoPxPs8JC0/PGt64PVu5sIM4WQ+HA6hj
QlQRusTCjds4aopwCcmiQXwNVbfcM5BpWHIA65Q8YY9e4a4npoWlbsEKzSEovL19
EmfiC+48akMADc8xJyoZ4HblcvhnoSDMORs2WEDbT5qDowkG0AKwCjsNUmPg8VDc
zDgW/Lu8mBR401cSZOsbu+AQD1zLFpRpp514MVkPJHj7mk7+LGFSYyy7HXzvsE8f
+gvXtzpel9m4Lxu+vDNKD99NgrxlHIyafIgqFUnE7suckhiOTouuEzCm1AIL8KTL
BpGQJy6j573NqTnmgwOJ9UxSQitIZsERuhamL0GMabHn/1twNVT3m4g27vNaHl2r
MhNMv08ROUs9MeDANhNfbphJMrMCWu4JTjMq5em4uRErSIEdWWCM58dN2DOrN3Qa
hivMXPM4+h6Bc6qAZvNZrR2UyT4kq3GgeG5UNdYkvMM6R5IPGs16XKQvom0X8Q09
YLqjBnCtlO5d+R9FHXqB+EZgaNYbVejkkBrtD+tlNv5Jdb13HnZ3pIG2GkCnbHY0
zNNiguAjyspr0fXYF4yUGqqHD2Wi+ctp5fzvAFjjrBQR1aglgHmQTYq0U3XoNHlQ
KwAgHCYtm3XsSuAr4gh8kuLxF+q98tb5wXZkZl6FTsoRWb/3A9P20ZTh6C9f4nlx
cHxSSJ8pqYBmhfrmBx33amrVWzEgmaOQDuSpbryVr3A+Dj4OtWDXpHhAXUPqgNls
OyTEQJPugLnQCZWAFoEQD0UvHsLn25QcizShH17y3eKH7DVYiJ0DnW1cnGEbUdQk
B/YRGMkRfk/oXT/DqNMlE+ChFwm/YHWYXSR/mVKeGDyzb2uHWHP+0npIAsoXCuGB
H/PKStIuhy59Lt/yJZnrOBfTOh2XSmALTVYl/NC8PLQCmaoVrrvLMZkVM2H5Pwsk
sfbLJURO1q/T+c8XXGGuvxkRknjihuWRSOMZnLpbYysTM7+ksK8WRNl+N/Jz2I58
9KBoCCiZJBIdn3wHPQmi7brYImaSC6IdwmUbm9Z6KcGBMJFeWa2kJ/IbL4AmQx5F
IshsflYJRq6TrbvMShvbtsb4GCzMNbpdnvnIVF2LpcRdxbGDtHWB1/Ad89Axy2qZ
/0MFVlUJbCVPtk7hdtU3aoZ6gAOFa/tpUWjFJmRh6F2EC66f6utTBTkUGzdZL2xd
cpL+Bota7+gl53lD//EIoSJ4g2NhAqKmaRuWskEIEc6iTJzNJT8osTGKw4dCGQWp
NI4v2B04UdhfUY2NtHzX1z08u0ZcT7cLiDKpv0ji/UToN0NvQGsyZDnXSsiosETF
LGgGajtIVqQUayCWHMCNUWgDkkYOADsi5iQ6SyNp0WGI5ZkSimL2JjyuwUp2vBKI
MEJ/y9+2H+eOxdep2LUfYHNCYa462HIu4CzfQHwbkPIdanCm6CHYSvZo7r9yU9qr
VGJbzR55f2s2yDE0eBWFBL0nmr09v8TZlrlM2YN4fOMCVod+WNpA4t46Z3U1C/sU
f1EHlAbTgn220CKreGRRMbXLzuS0lEEKzyoixuIIHfaTztccZ5IM7MZz1/mF0bZ4
14CX+EfqK+2v/aFxD8pmU6MFzxPxDqvOfHozpyXG4E0ATdMAhUCK1Zih/miPOXFS
+8zLjVcoYqFxz75Y0Ncv6kRa0KkFVj1zQUTWGkBVMrusABqyoIIfORbU0lBP6pBJ
cTBXxevasYQA8c2em8VEDtfIN+XXSmKsOxlW9KxJ7pGCDfogPwVaFQP19xDEwiCA
+CsVchIZq5V34/exnbaWdheix/iZx1yHW0IhivNNOmAGqPrSZLw43/CLm+Ml/2HW
JoJXGk4IBIpbpJplndEUg+VlmqkMAnXSwnUt0KEXjdZ6kkWz+h5GosC9CCm3JlFq
4v5Ifzbx9HZnPhCzvwTDhTAmbZyncjTeFAS1OSsuDt0G1eFCCYjnY1cqNE0s+m2Z
tRjTSnOumDpKiBNu9nR1FKifXYxeu1zBbaTgVtldxW4EK2w1fVMoNfeO67fDda4s
LNfzOcvGCK20/VXTyNuZ14Adm733TjvSCQahdsx3KY8AGoKg2SWG8/dWSXTIGmSJ
7+lgc8uEi3GH+stJpDupnLI3TCd9Bzi48kDhGdSWl30ir6PT+9K/Tx8ipGCR2RIw
xgUvqkyG3x2hxxvZ6BHnVE1yhkc6+h4/9y0JRBlGOCdd8IXM0npgizkM2j/UMqlj
5/krKF5LYbWqZUHqQ5E1OEKB4p9M3HXO2q2Oz9Oh5PmXSKwkceEWUxx+AbOTOgPt
BKiUbnok+klAHmfIgxb8ZT0GnHBd0lmZKw4RBb9WeDCDiGb14uvbexuzirgK8O/q
2hq/wS5CuQbjr3o/2OE++bvN7LumUotpzHdDauFfd89AW3WlAhtsKNIM+3D5aJIv
hzSXI0T+llZsi76d6w1dqmhsu/TVHRHWmZ6zEoagPNv24n0CW2/rf2+BHk9IwvzG
uYjNV4O3jHV97DGPzRx40CN85PSVOZGU4Zn3379Je9ce3dPRhp/ap22bpNFrFE4C
oaoNPfE5/0Im88ub+rGHDrSTPO1ChJ0PaS2bNh9BY8P21DR3b3IqWhS/UXGg487R
wMai7B78ZQ8hDcb5wkRho8etO+0VIaZZeLbcf3gHF2wL11OFriZT4009ZEXaAapF
yCrH+DV+ahmyiTedQtI+0UcvmtnG21hIcQeXsk/NE5Ze04g/Qa4IX2Z8nfKyrCCG
haP1ytMr/uNTfvamMyVe25j9dsuqXM5EuZZZf397VYKVuLKmncvWG2LQ+v+uQP93
`pragma protect end_protected
