// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:56 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
CFirrKRbu3Ley6kfEcQXgZnDVFCTwCAiP3J/5dXgcmhjg6SwSd8bms/is28yjlK4
0ovORmb7hxBL0G/LNkfqUPKaRubBQHsn0QrkvyNOo6PN3S4jGQF9lY9hCu3iXmoR
3T7G0ReUtRmNWPC+Cf7oIVb897olJS6bxcJSncAUY4I=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6032)
gbescb/n2sKj1vb92V8nImxG3mUEydszeFVuhFwzwdNsvTInk+XSzjTLm8LiPyq1
YXkINLYDgCH+BEOca0dlHMQ4Fg2yN7HwG/HWVJEbxPz+PHpSITQyNwABNEyXVHBT
QzjnEY+ZWL1G4Vhe4VVPVbTJW5UcH8BoCcJD3lFqmwgN0WcWPs5WQXlYWYx+IVwy
IgbrfXNj4QkcyrHZHMtxsfguyQRxuyZZn4GUAkMP2skBBG9wpUOSBZoAS7y3eU7E
kGalquERGSTYpa6eiBCnRwDOpJi/V1kd305RtB40wf6aFKhObAxk8yr2kcDzKZ/n
+SYFtQC87fxIqLdHMOKNpssci2P50B0JCdZZztjMbPkmcciOz8KYnmWkQ1od8mf/
r017OdJz5I7LjXQeHVgXeWZQtaFbizsMN/tZBh24N3M1fehYbsmoVhtqqP5nXsCS
t+E+Eu2ER4S157IH/mhnkzru/aAA8LMrM7vfM/Ld+sIjHhbchISueRwRamSYmX7x
MCJ48bG7uH6y9kllEuMAG4vSgogc+8qdHZ32h5GBggY3qqT4NeStXo+XHRqQ7Vs5
h6dAsDKzPKDHUNm4taJuGfJnKXu8uoGPzfZrhtV7rKPPPi8hW4Nro5xlN8HYB91d
114L2+tdCuJRnaJNFCtuzjCT4X8j5YpaGBPaZfNCi9X8U1VlcmI9HQi/P2uGZdEM
hQs6kC/GyRXCQGiUYBx2zcIWACrqaYpg6Y9HI7e3fN4bcw95E9XLj4//ZY9n1+CX
lpQ+VlYsK1ueRwDpaLW3+6NuTQKKsKetRXCYjkREoulZ7hG2LtHn17eoNK5HWlL7
l88i9o2eaNcYXWDzrEJH5rFn2vxl8dehA+Pg9fuRiHEEZKIABioIWrWTyJmsiKmF
6B++48l74lWVxNoWyExrykzqfMgfjTNJwrqGaDsaVtrHAvVELaerz4Iej48oEFcy
wY6059TE1b8aQh8G1UAeG1wmAmg+q0vPKgQzs7p+Fdf7SiTUo/0uoV0aRnrjoEjr
1hrmJCa5q3grNy1upJL1AaGU5/5NmSb33OJUBK/qBmqhvyDVyhDMZlnX9/wHMNXM
aNxVI04ktmzwtmotL3YKwJ9TySCjNhmzZpLv1WjsgZ1dYmP23+5DpHZpW8h589NC
S2TUtlievGSgtG4P2uyw4guQBZ5wr58IBM6B+VZaSZjbwfTjj6hYOpDHDa/xku1L
cEYXOGlo2QujWypjq7E5zwxrocrecg0QxxQU8WwjTk5/QFaZayep2B7nNE/qIOxo
WIpD3yZ5NnICbTGNYIG9FVpWC02JKTVZBXKlwifjDuKdXm1IpPskymQBywpF1kba
nVsfyG/GLV8kB0uMxPZFZxC10q5owV1Z5jPX7lTocB9XYrPr7evWf/utqueeRy7L
daNNHHPtCVM3w2bV3YBFc6e/mWslmIUpMnvi+LRFKTrtujnFW+p2zuvUY7/rmbW0
MbO5Yv0AGp+a0o6gACC9jjenLbyXdI/1g+fnhQNkrzoZbRm9g8bVMs1ZtHcBSelh
M/wvHBq+RJ+vsCEOFAs4H0pZPMhcPlQjU5SWPjXPIlTITiZW/x8L7UycYYL+rqKZ
T6onYHHXK42OKP/9Y8rBH7BmklMJkzGYYk5yrHz0BobeAI1Gjte9hGVdzbiGgg0D
DiINtmrYVASCD7HBNq5uCBA5QBAEf9bmMnSiFS7Gf1MReAMb1Uk4vS7Kpy3Sw5FN
/p+KXyuTdjVdqgyVyqpMsF1uBPkh0R2ULaFuo/1KRQbUCNzyn1lAqw72GJMbDyXJ
aurTpG4RMXaPgI4GM1ghPWCz8xUFTuvVnrvf+JhdijcjCnKpZ9M9dQ47O6VEx93n
ElmjHXz1fas+LavXZwmG4K831YP4CSZ2hCCMEMv59Np59v2iRIlTmkggmJKxzviF
zHGkSrWoAfxa8BGt+JwD267LZvAzH5g8EjyL4dQgm0bY0oBjVgiyQHt0b9HziH8T
SuWGGayG5MoyLzwLqvtcLFTD/k9RfWZ9FcUpEe5bTmVpzzuWrd3PhY8PlP7DBjEi
OGJxUd1j1F1j/h/UIJDmOJ1pYCbyXNrrW0xBfMsTPIZK3CFi/iSWFwz771jWLJ/X
npoWxYrOkqGwmgqfD9STr4mKhMQhPglf5Psq4bEB91Q0GmUfCYFqwWvMXbEKBMfb
tpCxcWobAwoy9uewKb+xEBAEIVidtwNwZeh+pqQQJm8oohFiaQgoX5zUAe055ii0
0Kc2jDr+hVC/mav2FDZ4gAqXb79K2Fw4sHqRI88a+jkUYZTV5rOaQmL8q1ZPzi8n
fBKQ+TVvpvERxTgpea+wtOWu0RI3I0KiZgK8CRRCtSnALMvMFdH1Hslui4gztcKg
hB9QqsClloJXi+1ehqBtHT4CMHl8VSiMGuB5AEJOg3Wh4RhMFEjFqZUjZXzVzfOL
WBC5tTq95M93O/TKCfOT5dVlQPHvv9GND7XjoqipeVBm3Z5qOpx+GHi1PfTUBUmo
GKCRNhuu7QAoexrVJIRi24lcJPC3lSbZ3IEoAGvWbBFYYAOERUkoExlmqQqnvn7q
IGw0wqyN/Zqp3UjeHROZxYL5WhxEHPORKukALhfhOioDEO5aiDIsO7P0ZAm92a4/
I+rIxSoiWQPi8RYqAFRYGKt1Sd/A8ixUtsvdyj+uaPrvFURvC+aEjTlF2P5G9m3V
cHdxZb35NsUrTAgmt7zqhhIIjwWGQBhC3I9IRlS82zMxePUzdp6PDPuW316hMU2m
kAWv1+GXDTNO3hjO9znY6cQIQ/qx0BwBE3f92nl7CltcR1YPjoGYMm87uBXA/Hw/
ROk3GUHLA6LgFWocP9t+iC6d5bLPG5ZXK8I+LTBKFXKcA/BAevTluVuqTwAYDoh3
MsaJRhlE+oX5HcCZT+1TdCgQu8LHV4SQwZ1J1MMlPGW7p8kcK6bDg5Z263/y3lRj
0uZXKBU2i6bzNGO6R2dgwMc9vd1JSyRiKtAIItbhKyTHWzOsbv8eKj9MDCBbYiiX
EUboi43lztwKRxazqvSrXTyauoIcNTNNOWF4cTzYH6EBaVN8E3Zyy3+Cf/EeTxP2
4CtilmzfSlXhueHC2TiKI9cX6gGJamqJQvxmBAB3C9lvj5OKfC5PegCeWVkr5r+h
/ipvYz5+pYd660MY4zFWdCgTATJ+f7G8N1xKYXG3ufi5353vbMRJy8Apr+gPbXa3
cJIEaVTA9mjH4JR1t84waugpDBRvCCVvo2Jj4DfJQkoyLieXZw0E7MwivqMgRYwh
JFytIOFwMXhcWkiBtl87uKrNn6H+LYv6XbzfliQSyrQINAb8mrNdGjTJQlChLFkX
yQ8zxpPHNe8DWdI/UWh7b22aoMKtdbQ3LPuGM4gFqWCfDQyA3thzcc895OaZubDv
qFh/bu8vyNOjywTZ3siJ0YR00NR3WuIlbdGHDCzv7euObCBK7HY86jU9QTlamN3Z
FaNuKv+uVo5wkZ4D22P2fp1vrpEMkHtsmt6YQg/IhU/3u2loYLM/7M+7vSnTGCZj
tRoPB55hez6ItA3BsE3dDUM9Ggnv0xJ39Jhy/fqoA3hajiqiXD+GrWNB12zV29xq
DO+hVo2TG325Ljtklfj9U4ONIM33hJEGK71xpmJWwynkqhswaJXf8X/5ssUhYZpo
AYKuY7R/TNwBAwVd8nIxScPpi1C/pnUT2M7q3gMdPPlm2Q6IjdC9qY5mdA7c2bOv
tez8ctnQw2d5hFd7Jbg7wvKrD6vm1PFJJP3ZNE7ubqDXoC4Vn9YW0H0JcQo9nO64
sCWARTSnqAKBqfbqpDIZRURlw2o6NrITn6FzlB5WfpW1sO7ZkOYyN38uBkdktWnt
jaxofBdtY8VXtT1OrSPkedC/z22hwDSJcSmP1D7q2Ah5DVL/TTna9UovLUjGeCRh
UkZTmuBarpdVz8Yx/AbdTQIzmFyrUuN39hSaeZKF3VQ10+2F8ZVNrKPzZ52AEIzy
8V07UJvbULGpRmGjDPVPKp9xjvXVRcunny6PpiLwUmQ1PNA1dWmdpUGdw75g5ryF
lCywYTUOM1/HXkeNFG29krvSUR5y2ZkK59YRSVp8F6Z0+O+MJiqxLxQzBUq0pxxp
BVOKjJIXcHXmu36d/aXpdAKY3UvASJnV//ObkXiItmRBaIlBF5VhnV4cuCw5IOIS
2h9IiykmPM503KxxDPU6eGHI4WiwLHOhbNlwh3BWmWamPIWkxUvAVtOmIX9aSoB9
DW8EifUdTwJtnMIwNr8icAx1MwgjyaB+COaYJ7229TiuAS5n85d7RFX2xTXjluWn
hbUWZ3ImJJNwhlDoiLBESfVb/3ZI2yxvvaYAQgjWeo9KOj+g2frXw82bfGmamUFl
bnFA+AF9jSOzT4Hb/9lKjPHLZaAQcumBX/bTr2Vr8XFQWzhkQ5zUMM1mTylYKLII
Vlpz+KiU5LMC2a3ydgfqY8coRAjtzCDMSuVub5EOVblu+L8ixcdW18v+Xl+CwTAh
wMzlN1YhNGYU0IekHajcZg5PYSMqeViO3eekjdihYYMjlVbJBQD1EqrlFN2R5GDz
8Kj54rHb5r2dDMVGSj1ySbsrmBDafSPzrdUUn1KUMlrxjI0eF8v4ZMvE3iU4XED4
vRiaPoO7F6TvA2yOT/WUPBkbwIV8ObQaTwe+FiNOXhZ1s+59PTi3OdjeT6LPGuBd
/3Kw8BrTsX9GVFAuycV1V8iNVT36DtAUweBFyZbTizLJiHQR/ES4iJGxzPsqjvD9
dULYMbLTfu7T6sGKxbaFd7hqx4qIhv2TRuTbwWkniXkCKJe8IWvA3xtdYytwtGJM
KZesRMBUk2KpqGj1+1zKBrExPxhS8iq/3QBR25YRp7r5ssfHgspXxyo4FlJ2ecrY
hVeiq7MlaLOvC5xfZbBgn6FseHVr7epjHGGP8pSTHh0lMVKJAmHqSrzIim1tJyqW
yYbEgKZposFKJ8/3fEGS1ZzZUAQ+vg7PiP+m5RJthvRoLVBvZImUtTWxqpikfKKH
QnJ7EamqEKONIHmVGr+iWtkMarU02AJljC8Qic7V/D3H0xFIpQeEkiYDthNAyjjR
wNOVfd2SrqblEcPYttDnIJL5cAOS33nrYOJRbPyPMGHQRaCqNrG8vdGfNfwd6fXp
JAqWYpREP2yypF0NIWThz3JV+eD22VWxkHxezVyNXHG/Yfj47s+jcmbA7L8dUNS1
H1EHICElIzxNaq/jCrYQGUaCvwOSjg8NEVsS7RIINtYYQOn6fwtxras0ZrEp4vcI
Yapz/7v/PVOlrCIaVKSl9UnPZIstRWn0/V3FsxfEnaLdWtP1V7BHgQbC7mcvgvTn
B3fxk0RdlsPsuFJPpnYwlsOPBMteKfJVX2OAcNRoIahBxjGl4HKVpqTDn6XU1+9h
imgVw8ouIT6Ea7+VFeZr9zY0qxlkvCdMYunSvLX6W2MjhYf9j6XLoa8wwxC33AbT
r5KiApsY48TzVwMMyr8zwnkclaTwU3YKhSgeav8Kvd14CEzeWxVCf2QmQg8MNMa3
ukxv1fojNK1kSaq41oN/2pXZKAvu8OupfOzqgLSSSuZp4J/jllEY64M6c/Or7Vuv
fklwURToiQioHJg7KgAZ3+I6p7qqvBAXIfB54IRFLrJuHe/QTKK2QmEInQgosEtO
tS+Wammlh1wQPLuyuh+D2scDb5cgXBx87QbB6dPloqZ6bv0lk28Ph2LaaXUaB39G
kSgjpNshL28D88+1eNalT7QXJmypNq2mPhez/tHoXNFZGd3bEZd8pZLApFRAmGrm
RQiEdWMrQk7fyWby8P9mhmBqT/ZjdUZw9GifyGAlJPGo6pSnzQjXs39Ax2VaCNdq
X+4MH2XLOHy0m2m2dAghdUi0fOi8eHX4n5N1FmaPoyefdP9yEkuWc4In98oTmj9K
yUIlKOvyducl8JPpnEz/poM/9UEEJVAgtHKy1A6VWMm2HUBLMC1UEzQuILNBoUTg
Vg/kWg3Pj1D+gKDAZKm+1888ZFN2CYwVw1jczUyPXFOpmkrg0UFRwks2Lwk50t44
Aa4VkKH7/3qeeMD6aifIebex6OrF4Br33ZIA+kDd/90ctdO7fljjy267r7otvUhG
Jj1rg8nCOletpNJpDNvks7EiYv0Wtce3Wt/YBNcm6hETFgwpHFk9/CjV9jtFSFcY
ubOPwaZAB44gCUtzLBuyAS/y0RCj1i885SuK4+iDxzkwVtAlfloqhJAhVjszGl9Z
sE7QS6vC/ikzXirtYs/IAM7RSRk/JN16C2iMv77S2R1RmwMQs9DgNi0AX9471sDR
bWS4eZX2pwFiDJgdvKQnNBqmXeo0JmL4gws9Huf5KUhdIqr9vWh+1xE0jD+iPYWZ
PgGhBBl/Rtj+MIH3sDZfnUPhsxRVlmIg5reEP3oVdacjG6BPpT8lKq/CKJjPMgEi
twnODH6NA+lKAd8kkQkQoJJmhFlgifj7mYfWIXPttJcdLuEQfxtrdav++SkKdg+h
xl/jdBXMuj2doJf6udbQZPW4W24EWbfzFETAvFZbPlSOJ0F8GkZyJLzP+B2b1FqZ
PzW/+ArDU31NfViVkSXBz5Ri4EESRI1DblRfPNrCI8Z8E63iHDZ/H+0+mxqt0xvh
kT8x6v2XRDp8R5AW9LczOz95ZDCdScGaO9kBRQT384K39pAJ6+PZ7NIzFJq58Vqj
8WeraU5n0Sd8+hhXoACyiO/QKi3odcay7hxJRcYoXC+fEF5iWG49iA95BRni69JH
QQwbcVSStCUlmvci0q3wV4LzzItQ7Tg862rBePHnu4GoIuFjpOZQac/8e9L3j4zE
jRxC1q0bsZU8HsBTMjQ+HeE1NW5rICvh0Ri8nHQxdBXzUlX0Ag/1+jAvEiLukyLn
268jZysV+fWEKv7V3Jp75vaGd1lESRyg8JmeYBRxYg4rpDnPv/ui6xlZmg7n4O0E
UaaItOn8oUmq+OQy3+Asjyi4QMoiD+NfFRpg23tZ/sd4/ZljzxhTwcGlJU/pJrCt
/xXKkxRe5UdonZsTbXb8ZUMe8VqyS0NNrsMEFmiWZNz6sB13TeqNfLxltl4nBtig
5TWWsxBFSiyFJy3dIJnIVLpuSQ7DVTcfQOiM9oHZ1RAxqgYvpLpy7otluAH7UJfz
TvxCFtadWPtXSeBDFVF/d7LM43fjjgWVgoq20ErE0Kz5VkaDAw7KH7sgDLdtAyK0
zT4/ofCdPFdIXm5wppk5VtO2YbMoSCaKEcJUY63RM+CmZCoEitAeblxjQsYuhQMy
zPJB5bM9CXATLNqCGu2VdnK1Yx8bQLU4HPsi7JKO3BHH9owHs1bsydnQDjWWaNav
0DPxP/dIbb3CrNsij/unRYENQVJln+geNxdTpv5C9Nm66mTWLOW5yl57scsqTxeL
HOxuitYyckoBS9NN0BzMwXqbxlxG8BRAg74mANVELDqMnmyGnmCVaJyfSesGgK3v
H8pgXETF4JW6Iu2euO/GLFvEluxJDjKuAY8hvlowswJJbtWcPcgx/bA6nk5YaF2l
dD3CEIcYluV2YU6sDPHdg4XRmjSHCjLAnNm2vhOOYYdQncp5COpoxooOhuT4BbHB
zC4utY7jQm7Ij032PLarQgbfUXXXNTPMsHNMpDbgEEbZXQPJUSilSucpay5KmJfY
+yJ/Oogbr3r4Ry8qw8QZFpY5RALgpk5IycHvBoS+aRoS1EFA8/UOPInNSacHWw+y
muanmnhuq7VS+r8CB42sQo46teekKUAfk23t+WEB3FEJHE4J4gRDWLm02JSL+6lV
rUhbu0URp601vEjavKEf95IBw/iKelEYrlyyMZ9/rpL/3nqtvMLgBnYzdXwSfv/k
p8QhYVtIg+8oaP21wf8cbC2poyBluDA9+lj1AddpbpYu5HfyJZD8DkrOBfMFOOnq
yDXW9LNBXJVGKp/RWKmAjbUYBPWVbyq4k50lnxhXd6uWs4CW4y5RtPi2Kx1PZKfM
ixNbEUhiB1gnGd+SWT4rw/hjcCnBqNMrcOfX6dlKNv4Rz0RGex8pzDlRAql7AzRF
jcPXdSP1PGYYvxK8bxqZfYUtC+i64rN5DyzkaRphgao=
`pragma protect end_protected
