// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:53 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
TBI5sJpIxjWr8biRmZSmEnL+F9BfTVf6RyH8fqJ40Ebg42UKgqpy6gfs4YfIBaDG
djX2XGYigYR7WwbVauhr+m01KiPogaDSCmWa9WRK/aZ0GCM2CUMmEO2EOqDrwdS4
pvybumgZrR+P8Sgh4Ftj+1u3acDbMmQXVcRRm6Ipzic=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3072)
NjJiKCjMWiXt4+QSboq9jz+RzO7D6fbI6Z1+u5futVcPx5uoXOC04GUdGTe8/cpB
IW0up2iRk0zZtAqjFFm5t9o4C8sO/WSLnChU1f2jLXdRMIw6xKPgmFD0O4C+Yow4
qvNKX/Kt/9gtgwNSKJ7u6LFogR2Yjl33/6DT2UHhbK+82OqazuNeI9G273E9PrTl
VHJHXin2xbGaAsCSLZHf0RCZPLfc5xV3NTblADcaNvrNTwmHrBTCp+gYeWLYXS1a
Jm88R2fskVmxQzgooakbJ9lQ/oGoUWCqYK/oxJHbRZC1EEBzdiVzIHXsCCwmvC7P
s77A/IxzogqH6RDiFl8BqsaePZIV8cfRecV8JGH5kwbtJDliAgjlQu4HS5PGbjhn
y4iHMbz2lGXP6DAwhmwkoxrWxh+5Nzdv7QdvLPvEtAS/rTDi1uZY/NvtW3Xlncz4
S6W+BcSKw9I0Scxe6t1/HfpdM0/GW5mKUwGqU+rOEUt9qd6qn5RDIAwZi+EfTCKm
LoBucGF4sVxCynJN/rfoJZ4Pip/CAJIc+UEdEOGF7IZlsHSp4PCOOvzRLPqXS5q5
taMXCWcdaxDdWDz8ALjqLuPO1xw3692+Mq+FmmYOaOP22Zh79RJvxarjcVtKnFLr
G1PEicuIteaVB4NwIFr7hur93GBf3gjvFUmasDBEP/4F431yfWVEFONBSceN8/Xy
cwJIDcH8TGTWaO2vGTmvuk5pdolcGeUNuWfpvjzotlHugEO47KhQ1BxplEbElGGZ
ERe3lPyDhAh4xgYuO72VM/fwfTr2M4yiMFsm7YuD5FTsfUI3tcXAfwlBDMybnlAl
3EccaIFHXujspYhhpgM3obA8muEfiXPoN/cGmy0IiiUGpQll6sWJpuqPImyD06Vd
fjjxgN1Qlt4H8JzZeWxga1B/Ur3mLqMBE/Ya9+W4tlkSjBm2IXZX/2vSRomOcsXn
/lWtS7b4a/mB0xf/vu3dFDWmKp1qlO3CozaY7ka8M7qnUusQfHRie9hzpycp9uF0
r6GIREUYyD0kkzBJkV9qTNGUHqkWHVCtxtuUxkuYtGkBss7ADEm9CPySa+rzUuNF
JLTmPfmdMCyEnmSYwBvkIIVyafskkrcFjI4Mzcyndwdwf57jDUUkbYkkIQiAIUWo
WgGAZHXPtBliWe1LlLw47Bhf0BpMlwkPwBhKdzPr5l25JjiiW0AOWx1CJGVkdpbf
gm2DBgKEsNUZfQQr4I4FFX3Lk1aJirdFsgaa0UuiO/S6aboAqC/JF9BCoxTiQ4Gi
O745En+7hlvji+BjKbCoREtjl4laWiUUWlyRxXm/8+afbiZ38biEPOU9kRygoGNm
Oudfl2+GeuV42BT2feFRDiv9ixrn86M/hCsDq9vDfIhwnTeqdvxePDdOQzEx6nVQ
uf25DDncQJnC9vf58GjWESEPmPo/bZVo44/yYAYypqRDerwG3EjT0/lA4J5UpAKC
8fftD+31qOOVABMs+hKC2T8CLzBySnivaYGqxbgH8G58qwX3u+Ea//DWbn9M45Oe
V6HizvPYy4Kl5uJe7TeTzYXOUfysndACwmbeAAOmGTJRBG2oQU3VZWHQS50cBluZ
E7B9h/7cIhhCqEp6Sv9B9knwfrzTHAmkx42rUAgBlWf4/qNfx1bLuWEXoDBth5Sa
vw5fle93WN/4L6hd80Wsa5qWWv5kPkU6WQC53i/ZWcbDxyyeFutm4WdG1DwOLapP
ukQkhQirDYYmE4mHDd04eDdndYuig5s1+hXj7I0d9K58qF3Tw77tEYwrAczB20wt
d0/pnb4yQIgbErTOdKWTvWWxPs9/QRmbsUtPaSfehIBrPgN7lxOB1SSjTkcjXDxn
fQHaq9WicpEHcdyZ8LNNNYqKkFcgZ+zy7OWXOMAm/2tEAlUywo0nKQ39k1HoeLGl
SHayQKAa9OEOQLDU5DYi+13ykjKmYs2B3Og230CjArN5+4pkjmR6cIgaC6fbl/kt
K35KRDb1tQmnYOWg5oBj7tNWmr80+rKWwThED9uNH8nS26JidtEbCK783DgLSu7E
eTaZEGYkjxTZ1eGDM7cf+D5gBePpXc5akAID7fSVE+pc0m0ZRwaxPumpiXdmDutk
aYgcaE2Sd6jfcTrbyopzs6G72Mn87yR4TO0Nn1sbTjz9cxcMXj1vzHb+qRWwthJF
31Yvzm4jSiTwD3fOEvXhzALtLLEHJO8hL6dCZv7dYb0PsujnmAQf3TEpuAVqlFtz
oFGy4CyCUy7w8u6xDmT/BIppmIn8DPK0x3TOWPdr7BcW0Zy5fpkBUM4z5SN53jPF
4Oe3nrW5VGotPGOTJK0DDbF2nWpkED2U80LsocEwgQPmo8OA+G8UP7lIT4+xsjYw
/oTYoKbv4U0W5kVFZofEgn2eV1yLkJIYJxcVyqUFQxg3QAatqRfa+eIDUPe4oYa3
ndyoQ+zrWwPnbqJ08IABXlkMOMf1vhzxcTNBCLfzJn0g6kZ9MNyixPFZK0DkNzF1
AEczFRMjstdV9t4uCDRn8KPiPb1XZkF8M8gdHkzl5HvT+PkcKHD8A7612tA4vvjh
nImQTAUN+zS9GL+XirS4piV1Au41VikGEo16jthlSM1DfutUCtlARqhnfxBkUTEt
eqGHBVPouwFWdeRkNIiLTKVu39D7qJFU495xq3rtbkKlc4C2tojJuJ6Ko214o6Z1
iS7jE4kdlXDryQBGuuId0IIb53IXf1wN/3nKrjGKq+aAm/iZoidQg+ApkdeQ+aiI
d7qirxHaJZ0tuEo0PokFFQI0EpetUpMvNouYS7+Kw8JvxRiJ8EyQI7cZhS/Ja4dd
mIzZKnj4yNmtojw9vnV6CCqP3sqtOZhaR2iurDYSiSQiWuuO7LLQEYlevlP4QuVS
OPdZEdd/Dqk0+vP7/TvqyRZaIZHVPlPKm8YLCyLS00OPVPw93Y9W2jWEQk66K/8+
bFmp8g1fJ3A5COaUA/u/ZmUy1ysikCCdRPtZKjBEy8Xg1J6+IobEdLCaSURQe8g+
ve8U5+2I+SeW36KOAmMqB22wiF1BF5UHwP27Gb6ClgEEcAioqBvJ3zxQ8I1Y4r44
AS+i6m8REyAoTJmQ2k0sfmf1IJVIXTNPXfpKLWpx9QbihulwchONZeOAQ6sDHVwZ
OM4NCRBOIwxsbV3TvxRhuiCbyWMOhXltf7AgOcUlzPOokExml8h82yvpeZDpc8fM
609elymhgTyMWu6VAQ2IN3+ZzK4nUhYpxH8tsfrlsvFgLGm8gyFP3meS9c85gxz9
XdsIk0pC5PKgrqZbIv8ur4GpCzbS9DEdI9UTdCwCl3s38EtivKXZTch+0xOMSBed
J6APCb6j2xCXJQfxy4YW9r5Bo1YgHh8O8kn6tO1LB30c7BCeqY2kVg8yTHXAuuSj
5Yfx9GMORxdQyh5fzhZblJGARDR4UxzWUNUu5XmB49JUQGtvut/124KaabWY17vC
a84XgDtC3XCXTFo0BzgeNH7EjWqbDpq7135FbizZOnKSI8HZ0/aMmyfzPJnQ6GTg
ntkUMHtqnVjvS6rq9Fytp0gQq4fXNRUoa5KtPPCOdZXtaoHFjeTh/6GdP5SKF5dB
U3zcNBt57fRKHQWZUf2YOqVmmIyEMcdg3Db+bESir/LF/FgIJ0IMy2KTiqyCYInz
IxCZhrAqbN3IZrl6qOb78UMLUCP9ideEb7+vOifpTz8op1/difr75FCXJGQZjT7X
o/hNxomNIGzeMbwBS8otPOIargmKtrOmlIm9HGjrwoRRhMyhXPE7WnAAuJWCWwtv
3yKTvKbTLNg2IOP3UDKz//nTVcDLRh6hSMwmfIHfPwmnlO1wEBjwpDGH5t2u6MmF
TfVWOj2AAbUU5G0J+6J8tz0Ui3EDL+uZIUpfcVjXQlhjyp25ErU4Uj6G0gVAitEj
pCO8yYOQAP4vgiDAh+DzNQrO/WS3WykuIFag7osWx0M8tknwZQzQmzJp+8tlC9JT
Sv1oD/6G7HXuEtIuqfXVzcXLpRhYlN4cM82D3jXNTVa2EnRMEeQg7gHkGfskU2KZ
JqfbkI8WQiYXNJLg86iKnQl3Q3BM1CJchIX2v/tTBUqJf/Wlq+vi6JPS69HTN9VY
`pragma protect end_protected
