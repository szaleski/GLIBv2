// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:46 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
GsgfYowc/hDURx2HX87BPr0xgm21buIPhS3t7DzzS+qTNdsfzMFqEVV/6KnPEKSa
TAqAOxL0g1PCB0t7ArwzZZc8In/tofqNlAaDZCd9eA7XBqqda37PhXg/sIp5y3bj
qf6RSnC9d9qGEwlII0oPUsXI7+RMmv5oAMSMQFNFnF8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 9472)
3z//zs41hvEQ7f1okcF5q44GvojY7wmtTZPlGTpMZYLHX+KMNv/hOxT9sSLJvT6Q
P3DcRAEz5HDvz52MbLvf6raS4L+vk431tLAcVyYmrhsBD1lPVoXmhBGlRa9xKdym
kXiTwCKQl4cnRG1KP/u8hdw+qI6PauboRvzCoN6iKd+BBQQg+jcuwh+sCSxxC/X4
+FaGf9r5nrKuwJhuuUY7ywEm/5Tp9xf4Wo9xUt7PI7eyLhua6GAs9dxOGhAy2Tfz
rDmRERSxA4BH7in+CbfAnyawY3vX7kAGutNyNyd43t03cwDOdYHnyNDkc6dzicQm
vWI63dxJuDKmjUAKcJ+lQSh7xm6nrtfRxkp1Nk/toZcaV4jjJpyPO46kjnwSyOXP
vr334dRqJdLqNw8g/xsA2IL/jrqufSlDTTVUSoJpHKdx6QAMNhm2CWLOUI7u13ZS
JsT97rQvYwk7rOGGewmg2bZBDHF76Qm3NnJDzcT78hz3fq1uUmbcZ0hy21SbxHV5
pm75nxJwTGScEVsrsoSNU/ubGd/gUSOUqnLz9xXKY7DNd9r8nrod00rniy3lHzSi
nTELYFITiIm3njhWJq+Yu9eBvuS/yTvw7FbsGCwOpi4ss8vYjArA96+ULJmW+nQC
mrZJtPWvwF34jovI9aVySzdsAr6XGsMPgDd9hp52lbr9LKw0PW9ApX1+Fgy8OUSe
Nxg5o8UZg8YIQvop3OzMk6Nokf9ia6AL1H6tcX8gYhJwWxV/+j74to1KBb13aNlC
PCFFuRu9eRgRmw2aq0YWeEfn3/7A5jWD2N1u1ImQUZPNsL7yyytzfyHXwhgJUqNt
AuhpBjUn70rJ/ic82jj2UzZYT3GT2gY8F8fSprhJrop7jAsp68w7Pq/Z5uqzMM9W
ZzJDJi5NHw9FNX/vWqFBZqdQ/3to23nTkf4+zf/5kS4n+S9NpUBOp1T9dT3FKr8h
crAfAuWjMJKdW1qIKJvc5dDbNklk8TD7OGcKZp5sN1cxNdhYGzPaY8gv9sNXPGq7
8t5DAoeMKzYX3oUfF80+mytei5s3ZAg+aopXlyLX6c1cyItjzEiDwoZaekgKso1a
HFjufqcENyPl4tuIxp7F7EJ8ojovlY/MoCGQj53um7HTl9v9rlhL7Qd17FngmsEx
wrUKmQ8X+1EwRV5FKyiVd+b9B1VPmo6h5kT/P7fDTCCOklPViujz0PHR4g6CPv3q
85QfByDjh2n+MFKrxM29BP31p/Hk6s3hi9z5wLCKL3ptbLoeBxJwjtOMSU/O84WQ
n9lbsH+XcddBTvwawb1VC06QQoEuw4N78QE/LWPxFyRbG1JT17EFFyn1LXtoHTLy
vpmkkTXtoNcHOYBmBDR/4issyTkYk069nHDpavTuxNx/kaMwzIoH/bmC5fPUKpkZ
KTYTY7O70QX+rCWLt4bMZ1acxhE+Ma3SVRslNoXFtI5VVJcUswReuO8SCdB0xi96
py4sq26acvlXIyHkPCD6uIg1IfbmU2smPO2Ez3xzPLbnJt4hcLXTb92Yzuf5NusZ
f1/AJnGV5xDJcW9wFmhDIUCPcszFgbpE+Y5dzwGkhCHM1LKzpaPcyhJQFZ7GAyGq
A8KXceVweGGQVQUDZdw5+CXkdqDZDlbnwYDHBvr7TzU93nUHWA4ZQTsReGT3FuOz
dnBMJTYBtV8O3To5vWfORTw0NiR0r1T0mgVQlNV4qwVbEv5k2i19u9t6AVuThFqH
otnwGujzSw/XjuOZOunaPUWsSJNBPDcKOr/DUiOGIv7s1J9F2HGnyYgXiHiGGp7+
3EkTzF5sgS8yoNCn+WWw9tMUGlEVBjVOotMKd6qt/iknYNvO+ez2Aa8x6xUr9c8v
xZFXaOuG50nXIbTBke10JQkOrudwvwDmPOY/V9sgO+i9HW9c7YzTeZs3HNebpWAH
ufa20l5qf5pzLmnRzCbH1JoSVjEWP+sdTA7H2flvYARyBKDnLBFlf+nArGgnyvYB
XO27LWeFsHlD4phQ0AlH674MOaaehs4C9vRn27SCssNfmraNutOig4CXihSg12o5
/pKZEXz/eXzeloco9xlgkdR7HANAxnv72lohLRPJnuF9C1Yszc0K/B6k12sfv05G
Ib9BjTic0zdMvUY/EgylaZTM1ZBxFfLdn6art/aDfd5dlW1ENL6zrepAy52jjUN6
gJFEPw1mzy80uXSLXQo2bnZOoagopHemVMm3O69k97Ld/Dcp1QLtVTWpv7VwtQBE
W4T86ImBP9rGaS/25sxtV+4idYEDOjsPPLp9eCLBu2dpmR718SmR7B8TTobYhmmn
nm5V0hUe4nzfqU98uOpVmet6i26Qs5NyTLElH/WLOx5zLJizideKPE7y1hsOXX+Z
NQZOjkOuAfR+N1XsVytVdABeHt7kkMmZL5mk46E6Wpo7g0C8lzYvVv+lzSkMVGpu
0AsDbHBdJo6RAsUtA15Rup3ocmueWQVHv+q860HQ/3kocdqUM4KAC5nykOUYtsHN
QSGq9+/QoG52iuzEotl0nUeDoZWwLYHBZpDm29nJJgdPk8RwpjwrMmqh/PCJFiGY
dax3UpvhvrSHK0gEISRKsLVIv4bZmkeTzYvp1PZ3QtJiN2HWn/lQzi1nvhjLQzfL
6RCsDCdED2mrhnyUtrmeAeI3J2KdQ8xzgF2IfguKbENEzzL7F3r+o92zpF/X3NJ2
fmzBjF3y6Z1qJ+UriDN65R8aAOyxjlZP10ja58YQRuqgjviWGZ//LoqCIdXjFQ4S
CWBR/d52u0TZw/vzWjezIk/pNufCv8IMZRRt9y6EXpF3/atPTlWbuQNaHgv3jAuK
ocSl9BqzxymygkSfH5r3quXxXhbolv9Lzm8R5sS3isHawsffsXHSCzv99OuKnWN8
8extRdtlBHN20QMYYQNN2RF1X/mCxC0mlWTiXsLIBsB51GvsPQYHcd8DcfyAP4xc
KIRkg/obsgL5eLzd1C21OEyOL+m8NM1Kp1flht7rkwm5aGCCMxnm8pvCESejxKKn
H8lHfB+m2i799GZiPRYag7SojhwQqAIyKHdbtzpyS8NPcYPzPuehQO1qYJJel0Zl
9gzEaqSqxDPVVyEX1ucobIS1pbG3Y60dCOU/eFY5gp3N717wmX3XkJwbU4dBt3i1
b20M3beP7Md85i4MR+nuHKAEHlAE1JjbsfZIWR1cHHPELN2X/v9nw0h/6pKMgUjp
QK40gewmdr+cfQw3HylmBWp1TC536wQiKqeiXefKszIMAVaYDeVFYivHGvYO+3M0
B1Or3Tms5pEMlLrXUWcqgXCSNdpEMb2YWHofLXkDHKxUZRkGcXYktPwv1i0W4a2a
wLstF7v3iVIrgmnZdns+r+cuMjKW5myr1mNdeBZeGk45ewhGHV4355h95psawXt0
LiF+BJW6i1QfqlHj2NqoWUSKDXOg0jwPjN/hVEFrDctpB0bkGMkqViMmR6gb/8WF
81W66vnxqOF34DKRbt9yHiH1HpXtye2iuCEKoTrf1WvlBMsAUxWREQcgwdGTfldl
3P5Vr0rU7ihRSqjiQFKpINMrBm7jBawNIwxZMtst8QXl91VftZ05bn5nMnp5yFTj
+XfvXx4ZxSTdHLkQ/JvdtWmOQ5PWtep0ikNgTJy3Z5ozmp+LT35iEW7pVRr5PIDQ
jWk1BspfOhNVY87xbrzP3Hy3dzQEDyb/+HZTTKL39FDwLAqghfmHljeVF7c+OSBO
vWjck9edhzTJeGj0Hd7unhAHLGOUJrX4zsYUSSbZsty+92+fjtlxuuM9fhVsdnjt
Css8YlvzJNLsIM9hD+iwoztmNTesoCBxgEPGkVfEUQm1BW5S/9ONYFTrqkKPxk5x
bWz0DwXHI0Qi8i13z5kdSiSJ86ArvGJXV9aYPGXFICh8EQ85vyZRDNuddRA9sYPZ
jEKx4lBFBfb7it8TI3uaHOU/NVjovtveQ+TzkUtGu/fK8o5cfCuteIZY7JVadgX4
FjxmpSejAvXvmAvGSeXH1QyTNUvNZzhp3DxYqNjo92bwPRzIRVBosCV70FwmbP5Y
rI4ciHwSM6mP2CKmHqFNQpdi8oP1R9nB/DBkY8DxTS2v5NpXs99IG3yGtFR5DhrF
XX7vzoYMEHjrbFW5jiOVj7tgY42c3gJVUOB/7iizY2EDk+DmmXhRhY+8ATGbcaQE
2w7V0Wu3HK0Ejcs4SMPbhCYKWtr65CnUXQU/gUNEv5X4mCySE3vVi0GiUXoIRmrw
v0/nIoYk6lx6LppsSyIR12HnJEAFv2zrl6cSnOA770NinuYbJT87VaYMGO4vfUJ3
kqbGW6uvnO9FwfBaS05/wf0pHyCmjOTtkOqXeNzIyDgswriBKbW3Hdp2/pCN98Xv
pJDJ3n+6TAK4xmxKYf4aa8H9lWbuOvPB4WLQyKv+7buk5JFlxeba80ZNohUFkSuv
hYj4I3kDEPWxqfwy3gT+NW3w7k5TCbVeKuaYX1FDgVX83edI5np3eJGMsgq2ZwGw
hX+x3jcH4JRluaR6J7WrjFmsclMnebJg19ejiKYFFHEUYrPuJnIIUTqiLh+aa1VY
s7P9q2Y5PvrZeRf+3mVLOslM8a3NhLvzNjr3JRMcKkeX680Sv89Aonm93BpLcD8T
wRO5+RJP4/mTvr6Iww9iGwSmYDms1ai67/HQTHjw2GW5xOu3KWBVtIG6oCTGI3zG
RpIvARagJAfqpDdP1LxmqTWCFpMJUeW7kLtJ3l9qobR4VpY5Qwl35MMeN1is9O66
fi+UBt0J7whMmugJ6bZP2Mli1GYEfF4Ml6lAINsainlj+I1Pgt6zxT8TxXIkqWaL
joqC5jwDAKdikdsQaJpEeW67coyEy/j19HMNhCPlw+3hmFMDg4m20enszajipAFi
TKSMDIlfOoOnQ3QTX/bBnC9UotbXsoDWOosOvA9zxbPx/055c1CLD8djS4U+zb1f
jSWpkv/j7x9yaEkW0fx0GG0JLGcbl0YL1ze4ptifN1noUlivIjOOyqCT+xWgZTbj
gpvHK40kXFjmxU5v9OlBf8CCknQs1ToPD5MB9BQ2ohxaM6DANTzkjz2wHF9kS0c8
fucVvqqvkpHXU7SzvtX2kdZCACRKHqnfry7t7W2ljhTuUJW19MJx+EqLoC9VSc+E
Z/2lQkGABhGkr6A31x78SC2s43SqpYKXp6obIlJDRfswH759zZE8sNlGicc3NM+q
QJe7ZUmKGY3jieQY6ak6TOp/iUyvzd9ZdaOB/Y8b26QY6CPpvIOM6Yf3Q36NIHVT
vSd+iuKND1ShlxptPmW6GeHG6RdplrozsuvZQtX0cTPz4gKWVsikWgPP1Ks4CmqF
/lyyeNEe3Yf4zqidVqzutARzgCzEoo/bjHAmvLd6vIhR1Lh0MwlSgz5Df4cOsl2t
o3yzLb6sXq+JO1aFI49kzxKvnHi9gAhRJl0cKFnK3ZNSnyZTeDQ3SIHn/LAvugd7
QsiBkB/huol1xAiXFb1wz2MBDmTGACmFanZtMPU769VO4N7V9J60dJc/paAK1Znc
/+/yAyV6bcnHLjy6fgOsZXXlitZZ9AW/IunY2XM0HnHNx7XqtVHRGPtGsuhZbpWn
mCtWEPfki4Z+KFj8Mhpk4ZWfzMs2BibzdzIxYPgMPcQIy7ctV1fKi6m2l0NKznLl
O9upBiDQ3r94dndsaTqytm73+4A+WjGF0dN3JraUNr6yl8DPd77+rp2ug3/Hgm7H
6YWP3kSxpGrtVTLSASeNmtt2+9/CG7hWAudcgHU6EpDK2iLir6GjZgTOV55fu7mE
Nyx6/inyxBI54sKAqUCf7h0tb+fbYdwV2Du5afNYrFhsh4Oo9RRytJ3qgEw6bObN
FNsYh+N3Ywl1fHf/4Tt6X8nXQ4u0Pyspl8nltQPVB6vA6IlkgQ1S6XNY6jymGiwP
8Etfq1gqILTC/JbmEwOwxgznQkpHCUctNi9iWDhlmEjhMgyR2Q1Uz2Q2JGYiKe3y
roPJhR2VeL2CnhJpLAcWHWjD7MKvp8jyQAtsGYCPhaA7xaNbmYpIFLolEY+1vtpO
5KeAc/GUCTLMA/JbwzdMAguGqXtkXDEn9wS8M7RRS7COMbSGqKTnMVBB+2BM5gBn
KBJvlGS2v1LIjueTnXvuaza8xSoBljOcLdXIgGq+wcM0BmRMlWUkQwlgyAaV8lhW
QODPHfo6VvZfyaQ7a19Yd/ySFh2PVGeWRHMvvnJUpGf6tijv6OU3+uyL9Ar1gcSd
kPAs/FwQPBbBtWAQbDSujxrIJFvLDZ0UbgU2vhBxE9HHJ0ZsCTN1C3NYRk07saoA
kL35uJX15dMUi8XB2F+Dah+q3FMzEpStTmqrITlujH0CXXd1aBjJrYZhopgKTg5x
lraID9xRpQmeVmT9gdMK7ctLUiCtDhM5PA0gILdUCVzufPzdLuV3l73KWMmpqiCc
kwdmEzc5ZnEQ4YBec3anZv4KD8OOr9BqK8kAsm7eELtGj17ylQHRRTf/hYR+HwGj
5Eb0oltH+nm6lWdInn/b1TY1kf2u3VEJEij97iR9xvZgSe5PVpldyG4Ie4uAn/EB
OwETTNYyPfAnRjQTcOjtMw7kOss2rIby9bpde3FlWGs3C4ZtuL8IFX3GrG6eYLKy
b0fW9pJo5zqZTqFbS3qz7cDu3E2S2YF9YSLVEWVhenRHXx8Iqgkv7/4arsHJpiLr
XIltZe9DThA0AskcFxpzbTG62y5f7mdiUqo6THhDBuM2ZDNPqXnlQOkkpY5bB2fv
pK4ZBUm1c1pQA8JfcJAUxnnJKyaNCdTYWF+wElXGMr8/RuD4QmeVgmKTRcr07VHv
wDvFARCUVUnsxMDfmvY4whgFA5cseeVSO8LIJmxTPQRPuMG2s4KHJVoza2zU3vSG
7HAVOgnjyWTFDzQP+jGG5Hj79xSqOKbq6mx/qY6fLGvqtrhTsoazWqd/aYUSn3A2
Ahpxg5q64DmFf+m6k7dpHmVjYVy82MUGu012efQMoC1GFaqu/sFJItxULrHBCImu
WXZMnp2xf06bckT4m2L/SETH2JizIO3RJS+84TPZewU60nLILrs/JOQuTjSzAn3v
Oagmf/EtrTL6QWAFEYkYxG5Fdob+afi6nXMMxhN2Xl9uV4SbpIS8wEgdWmUoHEiN
nN78WscjzWUVs0aEPpp5DCyd78RY8gmfGdshxZclP5M3ZairsV6abYgPPbQ3p+o0
1EkhoKKBhS5WWTIlXjxgcAUKpowD9Mq1wZNBB3PghaA02Q/i1NtA7miAbldwtn+2
HIXc5szh977OdYm0YvghvWW24YSksPZidgVYjeOE0zV4kTQyA6NfwpKNyd2SjoPl
Tl2/sjNNbTU7w7dw++qizhPGBoSjtmuVDHVs4WGOTEvqGMgWrWJ0DaRM1nORVz5h
JHAiHUsKTiiZEnDQ53/DzMccM7UXvela3sUTAfAeS9gx+i6YBe1XNBuXX8+nKO4C
OA9IeRtJqdBIqQx3LbhBciCRpcHWtcrJ+ibKvthdjKDjZgPDiHWN1zbrWHr+JhCt
Soo+syRMs3BOYw9VZlQ4dcEaR3/4bDx098Ts9TwGTha8+ZiNPdkpe9V9f0bBvg8O
Nf7I2h93jZ1h/mYdxX3wfysVGJROOo+MJYdY0sEkjqUBLUygce9Qo4G+NfKhU+sh
xAA+QW0NiPSathD0XMWe+q7KxNVDnIdb/HZL4TXXEX1dRZ1RDVVoG9caLM8kBsQf
02lviU+qeOOm/bJMiYrpTTZn2K04prrDNaHJIXn9xztIlod6muBz6pBL4lnGOTQb
TWNpJWDP3Q6qdqgvl3wFgl5q75mD7s8OJJ+l+MDMV7XaHGz5Inh9LGCf0XngTbgF
qnuQqWU5SJ2ckA/JPh6N50rMoIkS9l75oSC/UtuvriidDTayWtUHmTku4Mx9Ccrh
pRwFBTp2P7L2Vyt3MrsDJ1escfQdCqKI1ap7yOtaFCUXxD7qfvXeHUWjqRGFZx35
08qzVr1ZdK020L3krXONxYZ9NbDJQm9XNa45pu81CUREDAG/1MrTgImWnWesgde2
cqoFvd5lWX96RUxUaymFbtdCp1GWEpEowK59N/ge/Vn7JFJf2tkDOy/us5c1RNi7
u1MMPMFcxznv+780mqAYsaM8RuvhBQmfhOt2jOqpUPkg1LDhCPfT9hKqgaD8jVce
i4xAAiIMPptdcAUGYSPVWVmDBFjZucNGLn5+kPUEfnZQ5dVD1v8R7BAIpaE9dnsU
kB5daPHRNCUgTAE47niayWD91XIKBC9nkw6T5fS1I+8kO+qOmPwe+g1ouKhE2tnM
lsEiFCYneizceP+0WPbzbJRHnT774apSX70D6hLOzKnzLsaPy5bLhXcOIWeWZaDX
YkBW2UnqbHQuqurPa29ChUENQDuik6nHR00YXLU6DmDLG5hUVooYI+w29X8g+yYw
8ObnfmL7tyX9nKk44lBXR6mBoDwzJyfXrMy/tQstElpM2AvFgydQSzF+90MCSHcJ
YNbgNhwtl6vqu1kqR/SjHgvrsSaCbz7f5SspiH/FnEJF+beP/M5w8TjcAH67t/qE
JQs4Jy8JzE3kTRt4CZ/km5lWHQx9fDfYC6T1J5VROntPUafppIBWuaji7JhWZj57
HnahLBTmdzI7FcfpG2M+XRlhOkgtwLAE+VpkdUQ9bbnTyPzy5N1C7c5a3p9LpoHh
lHDxiFRX3egvk0V3gHdKqcS4CpVkTsrD9/9R0Bgf0LEyiuPeEqNAZBApu5fiDDKk
7l2WnEdl/TUeJzfDbBPIx0kpDNb8wgfG8WvUJkNGpq4GsZVypgEzopbGI2crL6O7
3mzVdeJygHhvaR6oaGoHHp1ZZcpg9w9gDbkDSM2E0LMtOl2vwBBC4GS8M9pvV3fy
gJ14PANBB5TNQK+7RgSEL++RZnoL8mdOuJqUe4yXKGtnkAUABnjkPr4oc+SQqmMx
IMgqgr8E6H5Enj4Iz+N4BiyU8+PcEdo9ANcgekhZLn8fpN7NZYkUNWs50akpgoG6
Jk2LSVdrKsQ7G7uEgR7dWf98U51o+pIqDI9afDGda4vr5UmmoFs3RTxabRDUI+n+
TEW0tPSQ8cex2Gn+IG9mEzhICvwogMDD3SBX5MdTbXq9g/UZYrvdYxvXM17gS6pE
KQx8B3QWyiIa47Pblw1pBIW0+9AK0FNbZ6XsPKT9/WWygDbNR8R+ZMjrlxp/1BzP
QAFVkjLWIvqwtQXFQcVQqEgt3yUkD+hygE9e8Acvayw0VH7EPTWrFSMd8emQywxh
UtZJFaVGVb1slezv9nVbJJHg0JjbhRnKikUh7nvFZy+s57JNqozAVaiTeXahpyLo
qC4YgNT6EFTFcsJ6ypr8u8egK4H5/dMJDmSQPTR2a1ao2hHcSoPVWvxipzhoj0Q+
LcKHun9FUnbqwZAOCYtlDxdBhk1a0GPYlZvPn/jQpZsbuZb1+13m8CB6Yh+PM2qs
oRWt5vKeDNigzs5fVEV8ODupYRX1JwIMCrcoxRi+JyqmQSzfscPmztftJb4F3s8c
NhcjsadS83of5ZOWXOKnDY1RG4al3jfxCYvsEMnT4sKF0z1zbOFjZiiwR9fSf5iR
T+rbwkNYkPy6ZlvhwsvIcH8aLwEesQBHJkkgF8E/UGajkvWs/eVakKXj84U+EqJg
Oxvo/X1Flgwuef9uKX2yvjkmLthAWix1vcOAf07P7wBu06M+56j8EKn2kb4GPnoP
OyhkFoE/TIdQUlFj3o1qydBxb+vRawtLIHHn49X5/Nfxj0z14a0jAMqum0FYD9/W
ix961rezDEb5dqYX90CifOp6PKEs0lnr3K3191bBsUbQgjkSgQBRyURBvnUDuJmS
+KVRfsZr5bpnFfq/raVmmjXtJinx7OwUzDZMrJmVFT943sq/GIOwqdEml6/GJ1Dq
JWFAfcGuAOF5P88yqjnmrfu7We60M+943no59KJtv4eOdPdbDC5Nwk4IpI1Di779
rCvtQaZe397IaKsEAJGxZQeDoFbX/Go6YUKghlAOzY3iljvtej3ti4W1YqEpTwlt
sCQ9FwXBevBKk8xkXtOzONzZrOuwd7M5gZwnzPwWmLIYVKwXZWzaieaw71tVbyny
Slw21BiRKrLfaStUlPF42Io04qASHVBVgly2AQECOFh3m4IjRfa5ChbSV7u7tU0c
LPdARCWEJTtDyAPJhSj+gKt9CPdKzcKI9bb/3ZMBOHco3gSHnLgboNxGZ2atJe4C
GyfzliprjVyAeeyFgqdUVr9IzHXTMPQglvmnAk5HyYz6+uCN/2H6xp6qS4O4frP+
nUpg/EwzIaiYHG4uUfBg+r5eENSI3xLLYgbYMTQS6gZvMmXhjL/7GSIMng3BaNs1
kNQ174e5qRGx06tQtBGTI0qMXUv46x83nDVp7NASwHnTqAnv9Ztpd4FrNhA5FUwS
jI/vHR8p1c0WXsSa4kfMtj6RRBaLOyokG4/rQEBdxDwe+D1uLvEeG4X4fK92rorB
CSvTwT4KSpmts5du4UscYC8mEM5rijhzImJ2IT2xSRxeZF2wpgP9NXTqmfFddmm4
IckcHTAhH2g6WoTUams7ryyZCy6m3epssiJIvNwn5N0IlfGT9mXK0y6k/ganUZZu
avbfHIL/qKOCuEtcoZtgx4h19aa4DEFVQNxZtbkTZLAeBxkh5bxHDb3HWvLxzPP+
XO9l4yVkHazlXy2uRlYMMYjO5TA4/LTft1iIKu14wkzwhGUgfp6T8QvYew4DsRAM
aDeL/3czfcEf2mZ9aefdR8ibn89ZP5YrGs1q4XXykAFZs9wb0aFTrBA78CUGjHmk
iiOgQTwA3MFMcBhewW2b//ZpfnmRDppmhmG5LBU+oWnlOrQhEsetYxUP0oisPrzP
mD5og6XIt/K058AXAazmtar1rbH9CRVwZe1pODZ6UxYpL5lKtKSfV1q7ZjT4XvYi
JRdwqRAoQvpPRpzbv/lzb4hPSQYqaKJdHQllpVRRivtm/2s6sV8hkLQpSqR+vwmt
hG1WIwsH25O3Bw+ao6mKa2Lvm9se6VbbCnHS6uoRu++ljWawX9lBfeoWY15+cJJf
t37GoXN/t0jY//u7ZyoyNshgeGkZ+11PFSJNfVN2Ml0mC/ZovL3MqnKYplBsMnCz
+0tbYIFFMBYH+hEZHsPk1YBFntlPDvEDBccAQi2ccojaUnEZMZX/FjM1ELnuZ11p
Z6jW4tcDPeTd/MBHFV2b2jX/RHkxGPx8wP94vlnHgRQPwH1Fdnw2pOoIErve/Elb
FvaSzvfPV3b+laai76rbuH0jcAOjcVgegzl3IGUCjoA5Y+7pTt1qnONTbnMjVyWN
pwNKOV5QlnP4jEV6bx49Ai0V35bcHqY0yacFOw22tzNrnCxiJLQksfzxaf/SW4ry
pZARzxs1fgGuK238CmwAQUHs7KJYkYbmG+ekYkWqPmfZB+RH62HEsjnDzwBcMwa8
s9pdcQPGGa67NIRP+bNbPfoqpM4+qlhNBSL2jml8H/ILwlQ1k3X4coST063lXUdS
e0oQozDRPYr+XQiEz8MuZ/a1FfOGG2LzV2il5nF5UtzTIDBKwkI6MBXv1mDFZYqY
onjwr/N2iRT4unnu/KbsPa2fpcjgRGcI6heHWoyxZq/m1GuB2B0A9Nqe90yNGWHj
8LYE+Gcf5Lu0flt4hMzpmRVT2ERkJjBwWr0MpErCkA0BR5sXX3Fhavwp7KGkXs+J
6woMuucSCEBlfTBM8Fq52+KRM9/lwYW02gmLwF+Hh1DGfUui6EtB44kKD5Iow9iJ
rcsvF522H1vKJXP6obHfuzDQoddUKvlWpdbkJ+hxwECpy7gARzBlBp86jEp6EiCo
c2YDRi7GAzj83ZgofdcK8OOGPgU55+iusDA0Yb4Tpak2lvgHQ78IxuB6Ltg9Pkj4
1/OEnD4CXhexqgn+xx/R5TRABazgpFthhrRkV0OV/DB5tUbhHRkvuavlz5PyO5jS
9vBOWR2Tu603Zgc5kAqD2DwrcvB6Cv7UkL6VSh2PLDYD0wGJIEXonG0N6zpXBnaD
gGTF0G/6ZQykux63YWmnvCypFKG8L/mHaKtlKrFtG68GkUCL0qu6UUp4mlV1hAb3
ynu1hjhtQ4zMiL+0NRHQzWVKmo1MrlPbZ5mc3ZC06LvpK1hfhsnmRaV6exb4Ligh
rZWkUKBv0WVU4fkT69ldDLzx0k69lhuWqA3O6xcI6FI6rV52WebCFZMJkxV6Nagu
/tvSZeSxNzZApGGgHV0qZo88iQL2RVNCuvydbaLN8bhiUEtqcYc05bLx/BqtYdRE
mIVHkACTPnckXIm5qVM6/XI2mk71sU42c1HIp7cgUNgtIlahm3ftem2I16hvUv4P
LyqZwzN/cYTobNmv+eDaaAMDQdBdI+7Vy65XWXJFRVeBvbsFLeBBLGMoTzJ4WVLK
Jl4cSy4KmSjZTui8s0wfApJA7dRmJ7d3fS896YDYeV1I1x5pUYkPr9CmM1ag0Mw3
DeorWLzQbCseRkdJgUQTviHPFPgdplGZHzkimXwsHRUNVXj2TMUf9+6zAKqJXUaZ
5+WLICcJpx3hUgATOj4+COraK8RNXGc5oo/7nX+9ktRCGoGbD6e3DA3Pa5bWxoyM
K5W+hIFDj1MWe2wYmU+cQQivzMbptxxD796QwjN+bx4uyA7dDM/q9g0+FQGmrIpv
/JVyhWippOPzEBVVedCamQ==
`pragma protect end_protected
