// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:51 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
lMYTHwCH7JiA9WDdHHt3UOSOEV20CIKKkf2EmSC7Y68SJVYDdXbKhzitbBuPHIPf
jr9VRrnI9JeZyTc3X3cHkEj2XtqBjalJ+AR74R956PGapy20/kmoDOAyhXbcn1+q
iygoxCsWzcoqT44OD1DUoXClTc3H0AV4fTm08eBQBP4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3920)
EusIdEHzqG1IY0l8qEHGJwWacCiTNfiOdBFE1jJ4ASgco3MEicewQrPu6I6SAKWs
br4n3gKV2ts4w8G/SdKKU1fL/2naCqzPPigMypokdyettkhtvkHauENEW8w6QXve
WdqBJtM8WVVofP9oUKR+eFsIlofVhh1LsaddD5mH5uBo5wu2ze/pdd1wddeqQODZ
8aiFtLeqfQRVMfM/+UHjlhtkSJ3H9YAMVe1HG/7nH8c/Nhk/l70yAPk1rwlJXMoY
QcwjMtkX4ZJ3X/XlTE/Js4rSO1om2m3VX9KZKX+rb5AyWf/9Z0K/4zIq2Wz6HA7x
+bQGoVvncp0/V6IkZTT9vbwJG+L4Fu1GyLkTS9tEIgSuprm+nYFtJ6a2gIX3iMQ0
1ti7wv2GeFuWRD6vonJQ1wT06ZeC93hN+YxJLNpWcAZTzevRNH6YcEtF06XXVjDZ
QexzKrXBY+31OtfgkWa7dU4a0rYKrKFs74xiZXJ9gVtTkufeLM8Jk7hEm20k6pJt
QB9VraUPptNYVNx54w2E9/J88J/NWMFPG62F3D+6TnbhUhCST5092hs1mAQIROSu
ckwBy/TkKGXZ5XE27u+KBvqk3UQs8vp5TBowjB6ru+xN4sja/qpFyBB9C0z3fzGf
X4nSCz7qwxDfibWgPp4sHeaiNAJ3o7K5O3HckN3A2T1SfTqwO0dBn9X6mHkELDFP
wGum9feUXXlM9FLNoP8OZ9tls649RPbIiNPggF0lnnrIJmDsUmzK1aUbKDa9NetQ
+mNdQs8yOiQRiQ47byCTG5hn5JWHEYWJywOBAxv25mKP931iulitw3qGI+EdDRYg
zmBjybBohMggg+nHkjLrqX7pE1msXALn4BaIwi7QGK9VpTkj4YSxrs8TKvXyPLBZ
OEr5/0PWMh3l2kwdL9cjy9swKLLDfsHAj+hvVzau6f1WIvXzrwdTmvpmSsRbnWSr
5ThQu35NBoU2sdugufJcLQJR9NynoDaDa1o4bpyR9Ml1WX7RaeXIz1zZgW5KPhT4
zNCv6QFynSMeaYehP2eIv7RmqY0SiPCvN3Slr0GrKWZ1ykQBQac7eInvehwsQ2/B
g/X+aY9p4jDsHLjerAKLsnF8ZTEI69EXT2u8GgFp0PIYeCvN582joeyy97CdHS89
2d5VJiWj1tAP6VgodFlhZIxgKUg8FBdVK3Wro+kUEL1lCNHKt6GQVfNHzr0SNWcC
HJD+anNvPO/8W+77z9bsj6mr8eOc2fZQBLV24LPT7TCtYs44I5+Ygej5X7jzBLeJ
JWGEkCY1DgkwFGJwhxY2Xtyr1TljjwAIi1Tx73u7G+GdqAL4y+OaP6LzgEXiKFPW
oeNoxD8GnM+TzsTcEeoVhQMaVIoLXUqHgAcNhZgv5PW8JZxUb4WRKtB/+9E2zOEl
foke3a1VP6JCb+w1mJBtR3V8oaUu6P+eqiizwfSYW5/xpjTkUOysc/eWNI2rGXqk
wFHGauBo+qZLshqjxtxIvlIOezFomfA4SjQtoRg7cpjP0KCE1gg3we1+pL2a4D1u
0eVWoIsHNv4qKjLhW5ntDG3KC3fu8f9FNdFDqnXw3N+gba3RWnXNpq1dNDQwR8eM
EgWetZANcyT/EEWqP+1qBTH8iN6V9f/MNMQtT679X9N7zozhF9Qwt/Uc5Yf/+Cdl
SzzYm9DbUreAeRzmsG2c8NiaiCaqCHWdVvdQX+S0iVn3S5Q98shDWbFxRgyo+efm
Lm5VwELEpGvP//qbwi3eF4eHyh7vjgDocXeLJmAQLv0x1ePj31zuClrqMJUzm/Nc
67MEsVJCICs7QqysL6jh11WeW86zEDhOk71Dy3HZuNcct7T6VegkoJ846yIzXoK9
k3DPAHb0cBM7DaPYHqeC3xomTHEpNVnpVkcb3tDEdm2aX4mABOARoUm1dM2yclJd
V5VGBkpxrhFNtKUUEfJGqiaKzVueLtt6w+V1p7n0nAVnlVUwh7I9oBQsZ3M/a0FL
S5f+HMrtuoxfN0ejYbKrNw8NWCmGlrNOv3JNftQ3LCkc061gTL4aUui3OhxvRQUh
sMebCfeX/tA18jzdA3i/3Vy9m7aZEUyn9B15f6+LxSKRonZaX7i8z2+23kIT+A61
+l3Dc7WFZD0y67W9JNUfTXTKyoU3pc5L2+aSkbP3LiaIjNkQ0BmFgYELzF0aDIEV
WOYj7iKeS4aRp6tk/fNhs2gBbGyoMd/xmClNy6c6Vz5sV/0R3WUQY5gexAUSIEw4
qFOeVgde+CtGse1ODXGD73IL0y3MGUe9pRN8EXyIxEhfOMq3gXeH9NNSZLc4yWnI
Ir14cvyr4sJNqxr7ANjoWlh3V5D9UxvMGGhgG+MglxxVS6DwLI+05Z8TMXUEz3q2
jxTVBk/JhDuJ1oU5iCGFyfIHxDpgII2q1IQOst4Xkhnsx2IftsIOeaiQ5lhsblM0
ox64CSzxBXJIg8GFSGvWPYlfXJYZ8iNS9rADd0tuJDkpKNS3XIbfvCgeqJj1+yb8
agf7S/LcnRdiivWQOq7vhSWLJr/PJYFp8H9fKK0R+TGcidGhljppNb9beUy5Arev
gx+V9Z1gwdtV6GHa1ZmRfM3NKG1GaqlR9F5rsnodShSfeiFdqU+aU+WbYYEkSpMU
HaAfWiqisRrV6sXIq0q9YP/vSzAkxm8n0jiGu7t3WJGoAM6Wzi9eK6bcDenYQlML
oLkfvfs3xX2wpgMzZXM9AD+CfdOef/dy/C9zv/IuRiaORZGz7y6t+TAh9waoq2L4
u5Ylk3zsU7psEI28t9NUPmV9IVkKlNdqAlcsYmoI8HtczUj0lmlL1f0uPCkxwtHI
qUJ1iPOhABBebck22Z+2iPg2X0ZnYUNkIbHTGCUeBiPDBplhAJogYXqox5+rrj25
npCjwdrpXwcyebCW0jm3ul42lEWKA02gCFsjGuxXSJB5yfL076d6zRNRYZZPXr1E
A3aTOp5GfRPwfq4JrIaMVBVSH0rlVbQRUU+uMOJm6i93z2KICTTC7fp8Si+97lvb
iG9F4VG5DeEyn+N/MThkN3NyDEwaRijPrCVXAoc+P3Xrg3m5kbhzozriG+BXTHXk
vdaILMKlmBztzB/QRbTBQG8j/y0lFFcGYYwwN+5ftVyLv9shMpngoDC3A4H/b6WC
QccxCxp0pAvIl+Y1rC1+5/tp0nrNVMwokt9QGQe0bJbBxzqXoQQq2jBsWWd0sN+w
ql2ItfKs7jDsh9Q3P7blUl9XHUhhdJchG6GV42G7a+NDja5B9xnHxih9Xybf+ZiL
k9Wguf8UjdzdDyYuUCbYbzfhMpOHjkG7iPSBb/xn8DqtV5f0n5904SxamAMhdR4i
3nGdMOXHP8BjsFIaEzE8Ghjwr+sjT5kNTeIpD7WdgDfynkjHMBZKSeL1F+XQ9guj
YixjE2KnIebSNEQVzzlbMWdRbHSiG9FYYYcXmTlyAGg9qMGZm3QRaH24CMoUzTPg
NuKDFKqtgXFbFzcei9mWrgiH0fk4cG68JFAZZYfZ5NhrIefQoj01EOjaHSO6KCwA
XgUdZ37RLFGZPvTu+SZuxj0Oir3p1Q3aXm27ukzf8JS86R/uq9h2Dq53OGeFUStf
0/WyqebwLLuQI+WY+6X24SDEE+xGWqr1RpUY4zRtaio7ZWQJms2ZTJHVMmHkPcz/
bvzq24R6HRIIgj+C8pRzT4r730LQHRtd3cBgQVhyfoSC+VQNuaFWo+YKTfTUlZK5
f1mrwI1uLx+8VEWC7hdRljPgwg4VVb9YkPaS0tNtQ/2vW/cNEabVk3zkiwUVk4LB
HwgNIUGyzJDTIrqUzmTQJs5j4pnlBawSf85hhGGNzLPYhto3++ZL3i2lmQSViJs6
HTZL8H++8Az4jRe1AUNgKBBs/s96tNTooP3pE9ASwENrDrzaKb3Rn724xaPEdoy2
6iNSszZ0FFdcbkQLEBLFeBdG8TWeQUEQCeTe7DTIffk98Q/ZV62J6wdkrc9MUN5R
qmVaVinPU77VCbZ6pAyqk1VftoL+vRUgOI0ShfQPmZRLot30mgar36wjQgRBdGj+
tpHHXEf6CyeLeA1GaAR7orZg6/Yi+/eEKhSm4n3E9+hUDUWVT4z8/qrzq0L5Ttch
0HWrruN5wyN/W0HHGe34ayDJLQzjcUClj/HMkQFHt/cUEWLjY/Bm5iVs6VHfI6t4
54+Zwpbd4PvXs2DnvPyp00coxFVZ4fnbNiK2S5inoTNZCSmZ2Z8q6G8ZbwhFMpSk
08n4Cnhsj8QYhTeFQ+ba6HDe0RNfTt8dnTi1X41OmIAhsx/+dx8eDArxAev+p7LH
bsJvSZuA5pCelBEF4i14E3WyXhO8EQn5wajdwaCOlDzgNhLNbakYkDhpZnwcUnTL
XHR2RKqzqqvZHdC/oS/bs+PT6LjGmvSNzU3lut5Ki7dhq9y6T+mByh4eN/n1wS2Z
Dmlt+NiQPtO8zl0LJRmF/lf/3fRKrWDYfmqNo0/HpzgCMq06MOq7d+gn/SdlWtkU
095Z0hHM8KJET97ZM6SgQBVlaxcC46AEie+w/c3dvJ5nogDPFjunlBL2ZkBukfKj
lMeIvgJ4AiNw0s9BcehpTnzs1B7cVNzJ0DEeH35QD5ZR39mGx3Fq3aNBa2awT4fS
ybKSzOrzdY1YikFIJe1/Z7ch+wgOA5dzmHjCdiqfDtltinIv8kLkuDDwtcAwiVZd
ahITbIymIadwgpMyaB29x3eNRgW6K4QmVOkhtKF4BsqBF1eO1dgKm23rtaqynNwW
LyiIroJ4q5Xb9c4jSVON2QJpied7eQHcO24UVCH42YNC8AorMfiycda2qdNp+Dvo
kdtz62qL4/MJJdlqLWn8c2+1aAKalnFmxEpbpxv8TeoVUvmBmbjkO3E49NvnB27y
lnM0p7Jld767S00N4xiJo7KitPq/8tXQD0/JyWurNWwgVOj95xhBN77eZWNOw8qi
0eh414OTWrUOPxevb6TNgBX5QlIyFVKX+z5rZLdYXmSNJmlIbFU+QMStZqVNp3k8
meKzY0AFRYOKDrwDG5OF7mgclcv/LHUu2LcI6pFPJ9REQIAA2XPIXToJP43I+djt
RfxgejvqwBQaHVk7EQhheVbOajAMZ3Noozg2ijYdmMfYRVsqkvAmC4pDH9mTHEUE
SaC2oXYlG5jcDYtJNRGDqIL8Iq3JWl2Pa8P7kXfjvgeyuSPWgFbQ9K5R0v89EM6K
gDh/VKVk3KuTYbGnLNn/rHSuC3Bk9qsRrsSVr56g1fE=
`pragma protect end_protected
