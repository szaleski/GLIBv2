// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:58 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
MpQgkwzzB+qVywSFjGR0r8R6AEe6HZRJsz5BHliiYmlW02eQnv8i8v7HImUrjasH
ucEt65lYbCI2+pb7JfrKTLgT1GSCFilw0kMLWwJLY9hGOek/NHvahjtTsusbJIXW
0soxRfa9JX3UI2RybDgS8auewVtBScI6c58aMoTKlkY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11920)
Yt1mOjiIzI+tb+hHFXAt4YLGhcZ+xyFZUXS167/OHuCecOdq1n9oTf916arhQpdz
r3TrOV+5Uoeplo+Jkl3XxKLGMCHuTWHmLt2Vw1Gr5q46brKkjROu/Zys07A1n7gl
L4h0dSq0iyKhadJ/YGLSUw9Yu/U8tUvl7LnbkNvpA7fxmNHpzhFQBxUFS5svfJ22
KsnNOpSXmNhGbsM5wAZ5MvlEsXCl3QRLGY1NyoI0A0v2UWRR6XAwoYBBU1sLYHFk
NAOnEU4/fPJZQpJOyGu1gx5u6s6uhyqd1JWt6R1DMRPQ288k2q/mpqlEBMAB8jXi
r9pL/806K/4yUxANdj27K9hVCaFL+S7xCMVC1CGvbZga4ILx8069Q+XAVnV6+7Jm
Wv4qgZX1yE+rRLG9Pz6emZxlmj5zTP/Jze7/25J2wDaFUO2Yw5SiWUBN/EmVxnef
xKgfFv90LuTmC/6O0Ag3+6Wul304IXlh6aj3AQSj6v3PdFGrtwlMch7kTnTse6xL
FQQkp5c8zNPiwpJgW7GGHHEq9tTaxhHPxXXRuzcQv010YKLWlIDM41g1tv5wHlYP
yvGWeASImsJ/S/aCtnd7MDneLS/OCU6d5+t0USMwaH1r3alPno7ZCuAMyClrMe4P
B6rnvsu1rKooFZjYe3mvgBxWYbcmcwPKviZUZ6qOgojEHERi96h8/pnpOfxoL5QO
iP5CtSZZ7i1zk+Y/rfyGXOn3CZrzW5b4gbPToATLai9HROSd6YhQirSkeB5RtowN
gGUqKiR3EwZsJ+rtnvr6It3SQhrUV8/2A5MsHEhJi+xTAtZW+/Vt0wJNJTaqnWbx
nHxizKYHenEwuIXybrcKvcgjhfTZ3AtFJ3RiDOumTmBH5ZvimZL9k5wL0zxB4MH/
Ei+VsOqDiYZgt7dfMxUEtduCP3VuerR7a67gTT5hMXK6l6pu3Da1096MXKXbyRgx
BD9iJDAyoEIxL0GOv8d4m6UetwqQXu8TpXD86OeXYPkSJgxjOFU8q5gm8jRYeUy/
lOcb7fbB2/3O3P49X2D4I4+IDC+ckKVXttNgyT4n5Jpwq/cv/sTeo1yEJ3x4NZTm
ZqRHuBPQw1Pwlydj1cD/MOOj0ZUqAxF5DzM8/8s4EtHt1tGU4xHSHN7jqkLg6Lfc
xX6HynVOnK0UcaV4T27WYLJhswEAas4g6nkySFQAvemiiD1zqyPgzYVsiXHt4gG8
cXMF9J2A94bK09xRC8War/eAjBqqtRkb1dzBS4cCb1mheidq67MBmdNqxzKIyVf2
nVg5qjQ/vfNIglCFhlRYSKVwK7NhMayU/2dRptFH2ePOpPP4KucXedpCqo1yI5cG
woH9zEnEoH6uURs4ZBL5J0uomkNdM3yMEWxBLNLosgC/HjUKUNa48J8Elfpn2ROG
KUzD5/ImzLOynRDH4NnCIm00B3n0NOeFAxo6GKPTOYwBrb4j7RtpDJg/f85mLYJy
zxAVQp5KAukbGE4bZkRRr0SrPG54gk4e8XnlUNp/2eQq+pXMm4yF+7PeCJ5NS/Jd
Y99LrkaP8/aRiS11jaTdkoEo+BnAwFuGJuQA9fUMLEjRg+8nwRLpsDaSW3tATedt
vb3Q6G6Jp0Z9cn6SG4ph3uiqNf/ahmW+KwaqpA65/E0Rl7ySh55vYo5kQ4TQgJ6m
etOBIdJEHwd1xbFA/GsIRVU//furwC8rVS7v2mKtecX88IEYj3fWhQH976BRRDhp
fhj+QoWgP860ujlj+fmJ7JOAKioPNCs79504MPcWlPRKA+2MDxb3+meBHJnpW/po
BvDZie4K4SGVBO2eYg7ZwWGIB0boRijzFXaVv09k4tkQqQuYX0jGE8fVpXWd1JD5
T604OP+mRL9XE14x64c3Rm37n9vj2v73nuvXtwFlLVK50JnEERocZEL7AinUfmTH
wkSKrOavda0cBj4KYNAyqOkGv5Lr5jYX3EKhAQq2HOGsRyT2rafP+b5TcWytoVIu
qyjCdVSTHKbxqwVeEIIqZp9+kY+LTjylpvtuZB9bZ0ccSRikilzJhZ7UBm66eYvP
znlELoWdWo0LeUAkirsT2F07wBw8xYu+AmZsog6SDKK9zqgDB5YmER75zu3KlF0s
wpCnJJVnQECvLjeae5zCaU1TYlaltBbfNZIB9DH8MLX2Zoa4kMu0JP5igE8T8jaF
/brV1WfMwStIv3rw9lIpY0CtSKHcK+0go0hVSCYj63BYWAjVdcGOHs9Per7QPeBZ
y5j1GdlOU/ByY3Z7qcWXVVQDJqr/8339H/teuxstERuMbPcHa9BdI975M1ho2xDg
Nakk32ZN7dQZj89fV3w/xG1vd4A94UII/ncnTnuOOGTqsDOdxwMvK/lBWSazgTk/
zxh8AQjc/NoRbGMGZ/9wXV7PLlZe84NQ1WLZtfugypKRIPm/3lgC5HHHvnREP5wb
/+qP9Yj4+4vZ/RAcW9u1NoVUGXeZWQ/esm6cg1eR9k+ivl8BnyS1LxEJx0WYozWm
F+K8Yq8+K3EDXihlDbwvhvVisKwdRO7BWzeGynICvjVrHVskTCrgWps7cSdiQH4M
AyRcCpayIatL8tUsio1ugVFPfXMR/AkAyKiqyVTcucIbq/Ane2MmEc0Voas0grsW
51Z8uGPb32TCkD5aziDTdo9XPIBYDB3a4tSkgzSWGCv8z7gwhx4cngwfx6U3j90q
oGRklU2BCGuHdHWI1fr0hIZO3df2h9yAOPTvQ6gT8Wviaeim/IHh7+tbJ2Y5MOn4
8WVVrRZvXU/rSNxghzKkqycuiPXNW5BBFQV6qpg+/Hhm+iTr2JYHmw8J4/KeuICn
0JIUtdiaNWXkhV+bl9JC6W8MQfThNT/XLxfDho0mV6BAZrmQ2zQo7VKRmBFYhorN
2BE0c4u+JtPzZA+957zrTw+PUg7+dKUJxGcswfF+uxwemdP+6kS6X8wcm+tujpro
DYI/kcpGi/zRAoZZjs0YHvNklzlGY4j+X+DlnadkfJlUCepNV0MumMIUq+QdqcTj
z+LNWEBx4Ujsm8yMQVjGvj4flXGqXTmMQIyQKt3r0FCStmsmBGv2jnl9z5Cphuj4
79mjmy8TRejei2aCe8gCTmOKUVOlhlF2xxDowv0anzNYezmP6S80mAj6P0slOY+Y
1K/YF92WTG7Z3Y2b/d9PqREtjY4/Uu3pDovYwyiKeFwKKuWJ8AfDlOop7eWlRk7j
ZU1vU8HwHTGo4ZOJ4MweEYOPEiZFW/ROGZBq2zKN3HhevWTy7ssKOtKf4geWD4Hf
UF6WHXjO8SqayyhX9nCoOyeAfLr8ViAfmFLTFGw3ChBbGA6B0pAWQa70GO0mCurn
sHUVNKfBPtbqANqXNuS/wkaPn4vewRABdWPpw6EZGzrkfBpQGbubrYuQoTPmykYj
XUHzhKFcA3nG++lYv1zgl3C9kKtL493rS9u80Gzng3d4SGVr2Lm7lruVlSMa4ENO
HAyINdKHCirWETp4BTNDP0ZvHmyXjRGgi6kAcIdk5+QYiGLiUSSa6JB0HJ1ez6WC
NkIGPFMKVxwWzt1AuNs0aCAdZvdHutl7aXxTH6CaDEeyocfsQg+hH7or10cqAxPp
R3xfOEk1AEWkERit2CqaObjdS/hJJ/C4Dfee8ZGKpsCgdgtK1QZtkq7gBuxHEIpu
y/Jm+4s0utpJcvHTvqv6T1ou2WQETQ8ax8wfP7WF4Hn4Kqml0k6U8v7/BluOA7iX
bar47zluaS/xwI1NKCcQmiSYbs50zz792x6kL342SENUMoFkI9J+URz8g5/efnKJ
gN+Hb4wLV528qiXYYFJPyEf8++EA71Ctme/xyaDG6Y7BVpXjCZAODNnVuecOwuxL
LHvsmlk2CutEeQywGqHw4cJ9fm0agsoxaqiHWZW5TFCVtszUwzBtD2GDSR0mYcks
BWSgKTZ+8pRwL5Rt1HHFpTyidLid5s1g7836w7nxVZ0yT24q+x8jm5jKQkrOU9Ty
kkg3mM2W03M30Wl3NeK/BC620VdAnmbuXucXEjBg7aNYcTBYuZE1ntZhAJW4QQ+p
16pJJfbviPzy1n8XTUvdKPHmdjNe+cJ1NaWbWrUUDl2xIOxrai47G0QDCHr1kE1z
fMkFlcEUfLLIdC6uUvPyTLfz4X/nXKLyiqI8vPNYX1mDsy9F3113R3hLcxlB7+7K
YrT5yo8SYrwuCYDNzyAR6Bws2ISLQ9sRItKqttsv6E11arIx4gVycKYOiRy3j2Fk
eWS3bO8ARZXlknYTc1FkyFnfCME/BM1flOALmQUECBfQ6MgWZVeqrh4Pl66GvvzQ
BIo5GKeG1DeTqYoZ3G/mMkJx7dGziLlbqgACdap3UBUHsVodWQiFY7zmqIF7G9It
pGaAbm1/7onpqO2/h2+Jh3XW5lQhnMMvPLXrlU5YhI1pdl4IvH9EX9RpFu4D/Mzx
fF3+eeLT8DHtYgBwLQPPjuIP6w6U0lsx6HgVOw5FNzC+YtgOuuGMbbLlf6042Ole
ZFWagsQQlVoAe+dIdzjNzMO5v824ZQ/vRg88ynKn7XTlb/PcHCFoW232k+nAl+Ap
Idp9QPFF2kFKVbLSaVLZR2e54uy25kyK/VW/nYUD2e6R3BKDXharWwlf+4y+w+1g
MWmglKW0egpIU2r9Sp7ylAWS+2/ReN5Lr1T5hLbPBB+QHMG5ST6kEG81NktSMJ8x
3meqIh+rYank1Zy8FEIsIkrljvGUMGXRzsbMHCqoqPWe0Q8nqozv+t+TH4TscZV6
Lly1DJ1IILvh/SDOktXx7mLZDhE/tK2fTxJyZOQNHygdSFlak/RytRPQpKrCD1yX
ejzsv8wnwzSPKLxqRwTA6FtfIYZHPwQVCGVI8wWhxZWtJE4Qe0a6Dy7vk5aJ8gXX
EMpXZCuLwJLj8JzTbgN6vK/51BUPsrGTUS2W47fB4tDow0wUP1/bRMY39pYRBwKA
MhPD6tztUXIcOCk8kL9fMcvEeCcmyYHZO1+c/ZCU0EoDOtbLzTlILRco4sBOSiW3
4LWZOUfS9l1zwpOJbJvpcu4Jw3YZSLDi379fqrqKwwYLyR2Ud7bDokJivqtpVVDZ
h6IlM/jlUjzgipK2vsP+2tZtSp19IT/6bIO/v/dwpXui9mDQBvrR5yKR7Lngj2Ym
rzsKCuZTtulclQU1BkNYymVqaAPbMHiE3nca6o82ud1O5f8sLK07HwzYLwFhUEJv
8BCPHd2csl4fJ5yu8IzZ78HsmZQRvL2JLCiVaLVwPauyxpGRmK1/YZFZAfFcQ79C
G5ZG/O6U/Cu7EOjWp2orbjdkMg/QkxAbANbBN72rQtLPnGJ2MAUQCKl44u8SBGbM
t253qSZidBnzIF+DX+ufg0kuktYCS0SLUt+x0ds6QBOID1p454sAdN8gx2r8n1Xt
uZM7pdb3FEvT2LeAbFRqW6NjXCS/I7hy/ez8fKRcBW8h46OcJNncWExjgpwSWyA3
bPGOy8IS0zChfaogqbKIebZ8KzVEYU877XLavMdZqa1pzvvsqkD+JfoqdwQXTd0k
H+SkNOjllIsorud1fm+7wb/xuAGcFk3LedcMju1BhEE9A3XhybRij1b1No6XQqag
yhDDzXe902kY7fgGrFVD0JLTg3fb/tNHLhXT1lUR63fxJAmIzhFP3NsEkzMjfEx5
+Ncj4CyfBHNOZYjyqGHVhe8mRbM8D/jQdCzaiWVFR+gLLvkkji4wF5QOWpxpUU6n
G5sHSC3N9k7EVXqrIpsaq28jf/wfNpjCbABnUGUQeLX4YYOIZj1u1/0fYGZmsO0X
JBfQh7KtZV8f9c+lsdRE8Z5iMcup4GRE4XkemaiVAib2dB5jXxOKT5kKj3dhvKeN
8lncdnjzLiEiDF0WlnAdrQPTLmahsyiKHYlcfcDWhKVOphBwSm4XYYhTJaTLijsK
HYf3sYv8tS6ZRKMw4lcj0jJseqt7LpEBHxSX75jqUHaTfa3DDlDD2D5YIFFLbwz1
1Z9V5ckFUBUQOKrqanj6xXWB4w/pERBUDy2ia9PMjFVaD8KXGMCdYmexC/9nJp4l
8TO0oFP1ZuSgKWZHEsNaijBhAAC0Jt8rM7mjWpBZ0YGbhBHRB72dEpE2cxtDK47s
yWNgAzWI21/CkGSMNFt+jBPcwg+9o37Fq3PgF2cNt+F+lkWTJaJaTaXMWrgnGZgG
ZRumYyA+PCPvvv9v1lvFd6EVEc3jm3vDw99Udxa84cqzIbA+ElIkqHsp5nMUo8Zg
5QYE5qOwygh6/0ucSicZlmTWXWoYA++ag9JRJpiE192E1EIhDtyAYP3TrJzJCLDj
3SbZI4bhtGQa06RwsalF9qxNp/cFheXx6+b69xNFO1A1Jms7coiCn2qQI+Vw4+yE
oOZxQzp8J8pTA0aqxOxZXcfQZj+MSWWNW1wMDh31VX29igRawTB15Rr2pC5Tt91x
L5FLALrj9LUOUZ9Kv22YOn/zj2sN5qSNKsEt2uVnoI9KivJOI+q5PafZ5OTCwSx3
SGdo8Zaa69G6ST/9h2s5niZ5CjmxCDmhYSAX7UdF15aBPfKOKpIdqrOoWg/8sDcy
ppS44W5kLQ3ZYzl+x1Lo1I0XUC9caG6WjKcuD5ePj2qoy+2MbDWNzs8Kq/Oey9hG
rtnLkZaeMKu7F41ftF7aJAbBdGn1Y5MQro9hTaUEs4wcwmNjH1WoEFSxIO7Sx408
Sp+ZPtkXICe60e71rUWd5vPy/WIVKaaZWGyxHVWFfjdA7VHs89uAW8Mr61pHELDt
B67SM8vHqnE7HTmZo/pQ5zwdmQ/jTD/dkbLpDjn9xJ8/ii8unFl7/4P6vRuh4LlT
WMYyUJSJndPAXZs4GQUPmICOr93taM26xxvdkGuFDkyeloIrLN8QiivX+KhZVIvu
suhWMhxiFi/qd0yuYwn/Wsq9H9Rap7q+TzX/tJ0WzMNQYkLOQQl4kyqKq2cWPzwG
f9/HLPXQz1PP3Fr2Ie33z/qYZYFFct/Xd8qSvmXMX8pFdpAuhn7RYHG50YbZNOJa
NEkOmMhLQTT/ITW9aKRYc7X0R6H+g29lglNKTQYjrMrM/+WtuzeWA83gqcahquIi
gTXvyNEgmmSjlBaLqykuzp1EFzpYcpNU4uh9+nId/y6icqvUkUX6R3SSQyA12con
/kkX4ohtdMf4J/k/A70SNl0i1APtb9yI2+yJjhYEsEjJEUqnBzfBVa6dMvyYdK4Z
OVp52prlbdsUK8bqSN4mjqWrRsg8Is/Uoq1CpPqW8Iyuf8XqGrJzRtewIxivB9o4
KlbaKhGQJjXBB1NznkuNQSPfZhkCWmUP1CSAEWrAFe+fzCIRGzcwbg3yLY4+qgUu
gq4NjESHcYa89k1yXewTlZsEM6xs0FTSTFxZQvgXLXu46/QlQvRN+yL6vYrDOv6V
H3/07+wH5xAa2b1H6K1c+KBhNxih9GKvWb5cSZpRjK9t1lYN2/xXHdNDMM1YQPsH
llfrSj5TAdkcmXMGIbS2tks4wfJ0nSaSxXCY63ZTu5HbJcnI/2Qq5ySjYOwd9QIf
fA7dsKKecPDfSKM1fNIVBJgj1K5jUeFzZJMlSjxi/FMXazC+2Ji6SWbgKfgEAZFL
oNB/siBkCIx+tuXdhyv53fxvofzv24BSYxBBAcjGFFTzkXK1QJNaoiCl+LQHpvdl
fPVfyHAuVYz9rrsggwbKVRKicpKGTZqwYi/W8uJvmwZWLoIeFw68yUOjbE3p5umA
SJetbz57cujixULuSdZVjZpcb2zEcYrkwTsj3bdkshv8HUv957xFMtvG4BQHn63W
FkqN0mmCpr2AB73j081cp63hcL5RsCI1Y/e90fSCj4n8/6NcXBvuSV+qcnObiIid
DVJZ2D1JaL782hSz5QiROvFLFOa+wPU112GuMct9jieJY8fgBLneGUbmHvWnbyHC
oOoQOkanil2d1o3aCFRuNfJ2WIppqfS4+yJBVuzeeYgTZ0g0RWTNfPBJ1dY4aytm
dPLugh5BeCbp6tzZMzIL4HEBK7NkODq4qL7IMqBZPnDHtbmot7Ald5PX51wZe06E
ZBIDZf71bSmB4pj/5342gfHBAk7s/l4Oo9FV/K+VIYnqmvxeeBUPd/T5Abl9IZfN
nLYXxE3xx/Nj/GUz1vBlZmjhSd8y6Cwn9SPcUQHkrIcZuissAaVAtJPaUrO127BW
rRBdTGbdMRTbsrAGgCje+NMyLmLX9QmGmlPmZ9W90CiEghSmSTM05DFCVzsBu9NE
YESVtGXMC6OJDNGT1eXwJIspUV0Yh2zc1qwXTBYLH/16Te8/IrOfViAmPmwpDJA/
PgvlFNCicNeh7IDHkdiLfFrEDlEKpPCQfxngdcKiJI0JLlDVPAV634k4xCD7ifgx
sKp3G8rpyJKfhxk6xmmllQT24GaB8WtRY20bgQ37OuYdUhm8Nt9Y+tne/z3s4wG4
riWzCImhJWXuEeLGlD4TaMLWYaFu+SyD2fIjzQlnKteYVtXsZQrWEdAk0tCGrFdQ
iu9+MkvotjQyD8yuxMNNqM9hNDhMFDYNO8HrRUnVp+3oy3XTI3OE4zsKmRdFm/9+
k5t1kPVJFrc/BY/7Y6L+0BZnURfLGP9Junk0DlvMgaULSaOQCIPEmmugUdb+9rE4
d0ywbv8pNlvXjYozaDqSiQQZD7DUXoqXXDU7s9/w94Moyq8u2SJuZu8gxEEcPUHF
Fb6aG2HKJ+cHgwyBwwzw15MygiOsxvNRdWmIWLdOnt/AzoHs/TDzdE5O7kj/em1Q
DBNf+AujUPYZMb/ZsPdFXtRi/08gpiTm4WqdmKlHIdwPufaa0qLh2vQyyK0TOpA0
SGhMmLQyyKOlpal3psVS22cjI23w+Nw7YLG+ovhiTc8WIRMSbU/3BDPdW45Hx/+6
or8jV5YEgt60rty3Hz9xHqN3YELau65ZSymvv9hMv+28VmIuGIdH7CecajdUhvRS
1jycOYbtGZT6V2WfHy9faeyvom6JqB5/wJLzfqrWn0E8LXaV4SQIa4xrmxyXX5SB
xvGMwqMCqH7dMvrdxCdO2rqGw+ARA2lvgqKq37Dk+iaGXlLU/nyjM0r5pbDi0e2s
dWxvpUJmOFFm9lMOuUAZokYSxQqv3Hh3ux9hAJiqq0L80CaVY16PsdB8Wklv+zej
B4Q44sSWoU/4p0Pfkpiks33SrxkC0/xFBw3M/PRQIVoHsqT7iLcQrzKvD0zcCxBp
X6ruWKX1ohazdVJ3LYje//Ge5wWsKseHDEulKN+jlTdzLrBgwxnj2uF2D9AJNLES
TyDvYGP94EQuhIa1wXt8sIO0BFsTfr+/sn616dgbFiqUFMhPLbviNtLqb+1AM+XH
G1tJhMYLF5kMWHPO1rAm1u7jRrZnzTtt/IeDtidAp3oOLeQOe28dpZ315U3vQnjZ
dJoLQ97pkA5ZsiM4Apj2uW7LAirARl3vLmvg8/HazJjqeT5859nelOQFCf9WUbXX
OZsjY2IUFEMMysw3gwMQxbxlb+GUhY7rZCqK0f9cEHZZwg6x+szYo8Xvn/GYgwUN
2tZ8WZ/gXXBz9K2toeo+XR23xYo6YhUf9dXOLLVzZRCgpMpjJ7Tlj7DN9HpfqtJ0
BFlT3nLc/G+u3YVgjSKpRNjSmYMGo87L1dh1xnAfKwaoRDl7YfaF2faOmlD4M32n
gStIfV57BHju7edlVZbLzWQXGioJ+qysp+SzDsVlXuHYOyTlJl95NcUFwQLN8BJE
t9kBiMZdi7B+jzwwQfflgMLcJ1xMfHloiSEwN00GvErW3zY9BzRUo+zzh+1FTQpd
Vs0ovhCsHisnWTGCumsZiKNMy2lvnNuPXxkhAIDBaOqCk9HYD9BzpfxerJpbgeDw
/WbySLXMALnbvqnJd6zzZ7AsfA1ar0LxAdWLE4bBzOQRUtiKmMwtYI8L0IUMLyfl
hR7lN46yLCQVwWDoULX42EiSHamJavXaZkj7HfeW7/eh/mzzi5DKdy7/fL/iweSm
IQylYsi8dv1LYwMdre6Ly4rDJFeHkgVMmv2ibx29HKwM1kxpwiwwxLpezncj+8Rd
XxVlyfDfXeZVrxh3H4ViocSV2LQBCXvlJ+7aVpF5z1EO0/ud2VAiG8AtYZj6nqPo
9Wu5ubTP5pB0pJeJ8aVmR5BMkIJZBts2iVVMngQxro4MWIJzRjcSR6d/EPgchLqt
zVpPZWagWn6WDF1dgZIfRWQcbb46gaWnCyDC0PUSBnjxxB4m9CDnhg3jgc1NB2rs
2urpFtbKsX3LJ5c+BByhwf8fRF56YEym8IBEIaKpF9WOyQwnoO++uRLIGqdX5m2Z
EOcFNXsScEG/FklGs98V+O1IJwHCvqIj9Cx3ragc4oeHyrDDvsNukqrjEB6gPQx/
S1wd2lxQQYAjucN6Ldnnzb4o+yxwkLhbKKraxSG9CAE81iufiN1STp1aa0TXbAgE
VxeTHilTxVCtlBjOKHH+z0m9xuyjl53M4QUFXxkeplyoyGWpUK9ezMBYbLUPEdtY
1H4BVw2pDtk548cU8luE2fAVdK7LyljAqM7ouu972GwJMvg8ArJkZLHrSN0cM1Wr
w3j7gJdyqpq3fhp3lUjcZlTLXYMhVNbrR43HDMDGv0Srfh43s8++2LTXGMh8rH5j
ZMErqcc3l3tMw5Pm/D0H/LmvvQcQSA3hq2hDcUJG8LWjbvpWOERuxIbrEgyk6lGT
zneijRFvdoTpiIKbdBtvFVrF6K4F9TbIDL1XNpLImfuHEXXxmmKCQ6K00Mch2QTZ
M11x5499Ik+T0tklxBn7tNh3k0fV45P28EMEfzyZw/qt5OCJsujUOxS6BbbGqDR1
RsU0aM3yEjSfJ+cf0OQsbiPetlpK6q12Osbh/chvy8v77CrFzLiRMnjp3MEzZBjp
6eFeSkhhQ8pXe6omoQobtgWuZlL9s2ZYzBCXh0ibSHXdrbk5xfaeE20bM8psbGEY
oxrUy+fg3T7C1Q+OyaQ3Kij8+uDkcvUVAs7JgnRzSKxZNCyalcaFxuum1kd0L5Wv
XWXV7JhGJiobH0w+uTFijIxuWX1NtIEz5Sy7smrPZLPQvJDfn1awavHvpJ9O8+9z
p+adMCZhoEtXdKErgtHMKDC1wblQL2Y1EkP7bzjQkq1tUwW4yxYmMogKXtEH6srm
FNtEDCYkmUaTWI70+ayH3Qv3WF7oJTNpLO8aLtN+ZqoV/cAJ5PVQFkPT2YQ8r3cZ
kZS9nh48+9HBBHocQOLdXiK8iqMAV0BfJ4TqJMRbhyjGmEwcpCHFa3W7myQMTVE1
NUXlWgO57J2PNtHdAjknNvb5pS0MqolyN6ihOeGENKf12mYAZJXJNp/zWVGt2Vyv
PdUb6L0MQb5Temg1fBIxZQvJv5ATSfovxWUmVTMSr2Cv87K5lDWN3uYWfBzSU4oz
d/20bCb/L6Opb410hidF3L9y40pq4x39O7sNCg6CFLwJMXPydpXOhG6NPaZdvxPc
XACo309hJFgGHQTEV3YPGTGGhzKG/AVsU5rjYO9zUNkZTCU1oDzn6DPLa6I18Tfj
C3mni148hnta5KmknoVc+s/wBSM3FpKbxox3sngT4Gvxb9BbFLEg1T41+7NUBa9g
cJmhBPX/m3qn1eFl0xLqMUb/CfO2DURujmSX5LvvdEM61vt3KGw43BL38FRtQFUG
6nRyh1+ZkZMsRT1EtkPKxugEEghc2WU5+dqxZPOZNYLu7Q7aAjZ9emsG5Ohghurz
sKNllQnpbEwD+7SeXhnCT+V93X7Ck39IzIU/CxBjVDjPWIR7TVJvSqQQurgGa/s2
TuUoJiWq6IN5pgSqXH88DRtWFzNhBYQEW1gdpLnzXzzNKEnHlyRNq3tL4YK9feVq
Yz09dETqT6njZuvcB2ASfRGoq6+YrK1HWGU4r9ZuuINcQ7uUSyZuJBAjzlBUvzO1
ebkmuaz7Ltg90uQo87Qdzj77m9gtSaxNUG5umWms5i45ecmTxwwT0JihMnNLz6W2
upomWmupFbz4gE3IUjUDVFFH/Y4Y01+dtc0MjR2XNL6dITYI3r+ceL9pgWbDhBkm
4aHKl3cCjyBIvLcc6XwwaQsaukYpKZai5gmGBX0ZhARVYobuzj/y+Cnx1raKDRYw
UHamedeJoIJV48KlfcZykIebdmIWgmeCpdTw4yIZghrxkYZeucL2QgKFTl4gwULv
Ul1wmhZ9JpEk6Sg00ArCDr2Aa5FvNhzPazmhj4TrjKIgNYh9ylGT2wBx0/g1Lc6z
I64TLbx+DiNGyePFfCSR1re40272GC1vLivISLgJxykmMhrzGvm0nxFrr4MwvL9Z
vligpCPHfJr4f1PN24ZqAf+vKbz5fpXgrX5u/v0PfD6Nr4L4r3yPU2xdXEgrUwWe
uJVov/EYVD6wLduwROUkI0zKQ92HwfdK5p1468Jmh0k/5T1eU+7LN92mWBWxoqiu
yHSIwxEqarGUF7JfneOucgpz9s5hEe/O3gkR0066hb9xJxU0ITTMAIFiBN83Ynck
wKyavCb1Ej4hKpUqknBEHVwPluqqII++fl1t6iIQFgob19iTpofCCZRnfPj+POy2
UnlS+ujQ0QSbOH+baXgZXCqNZRyUsSPg1ALxYns3azuW41DGwjyw8AE2VyZ5K7jx
Sfa6qRHinJT3zr31cNds/gOqkxEPQv9i5zIuk0D+qgeZKzO7jA4oMWhGsznqqoMf
V8AjrvCF9VtDjkQ3PbUbWok0+SELqPPGfCNu8kL9BhKA/uTd7+aoU66hRXpPUq3b
LP/azTUVQFSVa99Ukv7oAmCCjb9iGbHbmZkCQLF7+PgMiWHCYCZesHwGZ3MoRcAm
Pem4e2OOWuFwZVJF11nfUptkCmxUlO+Y1D5wgsqVMg7PP5un3J0TQzvAUITSOUaJ
jmLoElDrhYt9TPqhhW1mFqh1fO3ns4mT4u8wlfi6bjU088MQ+i3qDBM20Z58HUlp
VGMY+Vxy9PQyQoAJtolt7Cv67QBFp7kdxARs+yCDE64x8bFn+FOHD+bfLZadx7JM
zRzil+e5BKLZBQtMvqtqKdsQRhQcFjk04zYv6J8NGLXNL0hWBGh+hGGUXaFR57Wo
zgoINBRZbNW7kpGA91NLAWdEti19Yv2i15PPWkgluee4GWYfgclB3nqRQDer4oDh
al7+poZDviRPfOa7K6egx8pNn3Gs14CP6UP3cl2yc8ucJ6BkNJ7Ec4sq03pGGB2g
oqzFvrq0l7d4xFu2W2OmDUxxJYv/dZ+gYIjpy3GYGorTaC1hnbZtC12l5i4Rc2dr
YsGWY+Q1Rd4TBQUHTN2UpL7EmCdWCA01HGljGtK1MdHmbkyIspShSNqrAb8BS2pj
WSSxNyilEe/vgR1KEq17QYrXzRaz09sNvUqWdIcjAKGOAyWlKBacLusil3T+VBFr
/k3/oDzbSH74xlq/n78jruWUNunm1LYyp3yC1f6IdIHd2U4hvR+OyqNNqTmmUE4S
REvVPGOWdZnRUY//z7lH3W8Z6XRLdIwv4C7vz/GMwNbMv1P6kMyV0N142SrVBieZ
YAAu7BWHw6uby/0dNCVK3+o+vrYxb23ACPDqdseshK9SbwAy33bD7SIyyu0uxad7
XyYOtOuwoOgPrCpUmHtxic2cFfkQuF6cu0Oynqz6aI0lQdqPTEj/rTPRYrch6xid
4gwC5LztIaSVwur1WVl7w/dWVdH+1kiQoQDcBfE8I3RS0ZiXqcItJkiVgI5M+1q/
Pvt4xI8bYjh5hFXw8CzPijFhEtm+jW3kYJ3XFhh4hZiNaGaak+Cx0/Y5cR8X1Uv5
MpBtiXfq1z1Bkmq6tT9nVo+vWgbNiPnUvqd3GfMePWWugf7eX2YcbmPZqcccFK02
tgBHsGH9ke9GvmjG5mkODXy/BbLOunHQs59oNkdfCUuWuScWbNrmSAGdAl4+bf3l
2ECkho/aH2xpcE026y5GnnjGsmBsm1tgFMX6LdwtE3XPtgqf7F9aFUFXbl/IOIRA
DUfT+x8+ZbU0DXxjFdhXMFLntFEv9RkVBmvGrlpSDCJJhMelXXno/qk3PMotLIPg
CRjsBDyeMq8URIcRpNIjRGLIVyEwdHVJo03Mm2j5uGbv6Ogggl5qi5dgfLe5fZzX
CbNx/JrOeJNXHzc8ic/4ZnIj6maosksyIjfqrHq6nYFyZaXV77eebJ2QTEQprEnN
D1FuKosgZjam+IKP4fH/tyJR4dsGzIuFaHxFubZmx0nCErd8FA49lJ1rbH/mwoRA
fnvPCYp9c4EbGx1/IMezlQSsVPXrxYqxafkmh7NUcrjyVesMHzhJ8u/HUV8CxuOk
5Wg6x6/UiWADfjjIeCm9KMuQssRWSXFeXhVyUq75kysDUe8hq2XJgC8CEhaxhlA8
jA8itjN+AG04qTKjgMnL3+X9VqqL4qx3pCYDZuTXp9ruk9H8pc5UM6zqht4VCBtT
+DO42fcvYOpgcn659U7NbPb+RR/llp3fIitVQhDfbvUqqsoXu5WA7htfbvNe8Gwr
A8/o6QIzDgxcvPwVuD+oHVwTjWKO755yKGd9qS/lYsjmDrS14N+zfAxJjkzRK8zx
FjW/YchOaOdcRrr2fWbNE4fRlTb/h6ocyGUnYxUhxqdd//fcqrs25UAA8612v0TM
RSKdVNPvzFlh4cGrfpczsIWus3ond91kIXLW4o+jS7HvjWhJkudJxyv7S+2V1PjK
KyMJL/1G4l62UQpN4rXecH5PXbRr/BONGI+szweGGidqtKr4d20i8DitdbeUMbqu
3OizVZD8OTz1ALGhm0qm+w/DWA/cS9T3KGRncLNAD54JjoIJgdSOhsSvKmJC+YmY
XZDey+7v86RipE187XDk2/VBd8tgrWsQ6aEqr/MEtuTV9YIsrbAfGMjIsb/8JL4B
eqai31LHgrT0Adn+vceMmjJ8OJYR+Z2Ud3btNL5nAI06wUvk+RSVXJVgHaGAgaQ7
58/NV/mYpt+QP/o0bLXcr6C5L3KPQu2YTR1Ck4ZUpGfRR3QBHg94pEMfGT1nqS47
Kf0tO7AUW0IYZmpLdzZp40Zjz9KaKzLK0Prb3i727zsXYWTZCr7WduuyhiVXg5C3
QOK6OXK6abHSVqt93kgeJbe3dFvqVPZGyKkKgaCag9ACClCHhwAr1pc4UlYqzwcr
XfUenV82dt6Ew3z/Y5cCggWiLSicKD21vx5LhD+jSQgecQtMW/Q4pn2NJR4DRt9Q
oinomg0bsZcwGVHO0ieyUO/Yw8SKnAxBCInLC9g59R++29QN/KQWbN2DilYh7eg1
xX3ir98Q5I6Z9QYAYYFDCV+yKNySjR4bFH4TLB8F/QC/aoccCQOP1ktFNUiuEw62
rZD26Ri5qPUygzviYGOGl2TH+cP2zS2FsJm0825wlcb7gAXhGo4e51CkEHmUy38X
FMR0j3dXf+CoxhMFsXP45nWRz+FabJ5P3yPm2sthA0yKh3H+1xcJcZlibcKDkU02
D6ZWDiCBpT9sNw96jk5/peSMcif17ozJG/9/d+mnzIOBUUoez+y7h13rdFkPRleD
wzqxjcNLhKw/caBrwARTDpreYujgWENBkO4n7bcIAxc/uewNSAMZQqLn0tZDH1Tk
lhM+Mphai22UTIEgGOdbncfXUFdYbPLfoKy/MvJrVQbgorYfgHdq2dAjd3ruHXbf
YQiprKgyPvR7sANVbXxbxZPuLfCE9Tce9i3oQSgySV11AHC5eoVIU55lipLWx4fT
DwccHV2EYoP9HCqjVZ/2tIiU5YH5FP+mBUdhZoXUNr29c/v3Sff2OjtjRqsZUOiz
3qRkY0XmLqgFedd/aBpnZRbesFMab9OgLtiOEDfv1uUpdjEM1vOgbE9MkCp5tLQB
yWKiWLcBl/O0C7/1iICFWzHXCK+rwOxjAJN0GbnbsZ3kAQqXjs5ABrfQO8/rcXi6
OoIyX8J9hJpaLv1ZsLkfwtyD/9BUeuq8EuPGI4togmVzX7owPk8VlYBz8cZF1ddk
cW4ctaxyohzcG5u6m5W3ow==
`pragma protect end_protected
