// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:57 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
e1uuDizrAeXjXqVDg5MAwoatZ93DgoDVarTzkh2rfjbX5yBDO3K7sBIRytFGjHs+
WWrgtPuc2lzDNjeE26TNSt/VxFuDSDdVHKX6iXsmJKGw44CBn/Cem0k2D1tNjHW9
3SSFQcjNq30KVugdSh1DZLbnWhe4weEWaGN2dUY90Do=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3968)
H66cYU+N/GDuNeBi3VH0j0lVqvW2WOHAYPHhM/pFWUIvrMzzPN9CU+3aJ/+WlsGS
1befsY7MamtS6xB1h0p10Gr/JdT0L4gBS+FjgJvIuEIW48b/RtXvov+jM+2sTMLi
sohTR0mjYa5ZAh1JMFA5Ejw78LtHxNXdYxr9iJew+fI6EqXKfCg+f7IOz6jFStQH
w74h1roYBlj07PKS6r8X5HW47wUvJ0cNWY8HCsKL34Hb+pYg2WuWIa8lBVHRi+gH
NIUz4aafsQrvYi5gC2tF2XrX+W0tzM8YHsXu7me/LbS9ycmJLfyr5+/sB5BZ5lDW
Mdew1i5PGWFEPu/ni95EVjEWFcRl8pMNlTh3aAdqpuhRk8V3rcWXj8ZF2hDCIHh/
nRRhMw4uGhxsIMtMxcrWqhid8JHrVsyJFyonIFEOtL8heEqRz22b4X47H0Y5lSQt
htDqdsbisHKiXdb5WA/K/aRo8ZLM7tyTJMyDe78lnXyyct+eRaWEzjFDF6lbMFSS
Nd7GOqRyijI7mBJ209Nq87PKz7jeC6ZH07pwomjmEDclS/Mzj1yuPe5RUHh0nbpX
uI19MstPiYYLxHW/bCrKVk75ZfsHCIXCSJdwEwEkw9/TZnJS+MAfYrl8e/yIhnAD
/6ErkEDQhkxvTIzeQRyqlpi2YPgppM/iYATrtSFjP66fHz7aDMOcULVHhaB1QZYn
U7oIpFTc9cfCEuHx3CY0LZUr5C3VXyMCJ9vIS5uRLFpvfaLtlP38kMVstZkotVGo
p6vgynVlPk1FdVyYikBK0VttvIIrsr7bMwkC+E3sovCqroaXgGQuof5YOwyZwa5h
u9Jrw67bbLnwk3VEEYKuL2nDwQzpEksl5j1MdM9yT4qomwRkPkkx0rSNQnJkAe72
rhi1Z6Fo6j9uw4AMymgqsc6RW6NaGO98TKpSUgD77cmdb2VyE1zM+XuSpVXMMv9Y
lJgBDLzEhKdduC7lRX9z87Zv9gsJUDwKK0NL6zSmrVwfcKL6huspRYTUeVDKg/To
N4H+7YOKuEHsMifR4qnN/JDjS2NCxx5WyOQnbzeW+8kBJqNR5zA8vfAufPkS0HNW
hoRh5igJG+9/6cjx5Vc3uMLfwTNm5UIX89+KDvWzJSanRxmGTwBIQx1jP6wxLa8E
MBh1aNL533jJTOeXUarFz2uiKe6B2Zq06YNlf+6JZb2y5FBBkG3X6XqFEVQqAFGk
XaihWP9uDYIv1JIH3/oeMOzHxRuDtKRcdLCr/aqGs1HD0ecMxtSDiNI+GLdSxXqM
p5UdO8CUrDJ/sgjeqlc0acpR0s3mt+ANxdQWqjYXi6S8CiLCxYFee5xHDWB5UHAl
/s2BuvT5jsefIC6246wIrI5IcSpVrWdDKhNtohy/Qb/Q0E5gxqDun2eWCjqmsZoq
snjKoKuqlNNgvxlfuuoCgFOrRiNvWxPaq/nr4g1CigcnFX6lMpWKoB8ixPoXRgJk
d9mtpXJt9AjFO26NGHeLuzybA5Ae4Z2jxl3qBSH6gvYw3xCu9Rcuu+qE48LWZBsE
83RVJutFCCugRBIZve9kzHrtgGkrpfW3n8pvk+hkeKnKNHH1RvA9KKYlD0RItC8i
sXkIuYesT7uo4is+DfuIakvTceHpYlTmVez/J4JcmRziGOwKWwHU/2Lk7UptzHwu
zEuZ0tf+ImAeIC+s+6aJmk6OCPmf3efp3xS8ksmRO1Wk9iYglvEhwOgRoKvN3Gy8
vaxd0lPaY3iY7OyPhl287upiskuXKfkuuyV9majmwL5NjMsuDOJhTGf+iTBFH9xL
7IMpBhWMC7jUfMz9k9yUYsjOED+3UTTtPnVUPdHVR5fgOI3EcjRn+hWsYOneaL1K
BDmDJaEWf1F1PaS9G+1IYViFPvRRWP9MlTpnciXZXTUaIKtYAgWg3yID/d7FUxvW
kVAJUn3UeR5Yz6d+Ee2N0pPXOkwDomZ50LwrH+EEgjkgEykL7qwIsfPdLDKLlcc2
dSzhckHTY8An8iE30DlOXmIPkzIspnZhwSb+HsFsd/jt+T3Q7SwCFQHXnZQRKtZ5
LXwucdJ5Fjx4G9pY/Oe6XQA0W61lTs397VYvOjkI8WtZQ9N4aGJrgxubCMlWlFtq
mxYi0aAI6fAA37kn/cxvsUja5eKoClmkQa1u+t/Q6JZn5znv5RuZ3+S2akHrzBLG
nL7Y/ZNQWbvCsZArML7jR1Oefn9pWUUEVMjKK+3I/q2js1ZMjQ2jgkmPOXL6OR6x
tyOYxSBQTGo0e/d4S34FXjbb5epxyEeZ+8/CMRz7NIYGgYd2qDuG69fBpJw7vbIr
q2ayqDPMv6CyjITfXhWg1RzVLzHXBhAVH9+vcNCm56wBOCft10p5xvVytDNtyUU6
2YqDiEAfXtByWRq/nVMyNv8IeRsb7yi+FkLiFIbaowG+f/ocURgPoUf2oGvgGsL/
O3IGyAa7ifn5khmqjjjI1818wGXcQqGgRouhJ/RQ9LBs7I7XVIhbO8gs8qMYu2AT
goDzhAlK1jfwjazMGF12FXDSZsHSy4lk7heiGVPva55DBtWed0T8tNIYmmmiuCke
g5X95IfBwXi5uIa6hDaAZts9ReddL/ngo9L/KFEx3ZX0KS2Ew2Bc6+w5t4FZbKdO
pXd2RxfBlE9bOkODORkyFj3dZ1VUdW9DeHdq5SVI0a6HHH4+qrq5V32OYMnsFpxb
NFD80wsW+0MwQeJZiipK6BaHvOx7vP2ryTT/PpozUacLRk/7t9Iq942Pfzjz94gW
YOCYprHEV5Ixts5LVdGuwzOB1Y+uyDZfQmyFsS1PRD7drZAoAw5+OzFyp5zIAlDa
z55PH9kPlmI710uKaXPYYiVGumO1fRy/SOOV0ai9G9pc7P+Sf6zQrwW6Nso32oJD
K/kY2uxbbpzCum+h234L6n4JOLtzw0GPFn6foHE2dCn1VJOig70C0okZOMvmQ/Mk
hAgjw8Z+Xr/HVfBwXnTjEdZeEK8I/sCIBCbxJUiHsExe+XzBW5axFsfbyAuSSKUy
Y6L3T2mng0uelcJ1KbfD01phbsD6CUUZ4ZfDX0PS67Iw7ZXIfCfuOqDtzgRbkhyT
iPhbLRs03DN1WveXOborw8deSHKy/8sTIpx5d2/0LtxLDd4Jqx6cKVsEDgQRCsSi
Yf/OlMh7o2AGaQk14SGg+pSXTezUn9oXeKbHzn+dKN/+MnEFmzoEYhACoWy0njdT
1VYzJMoxW73W0VOHr1pK5BtL7GCz3Mhxc3wAKTgDYAe5FSMgYu2rbPsaleG44b42
eIM8msPPYiKxPgHkBvEM5Hvtn++SdStOfvkS9myk+VsyENefmACF8AFuFz6Oh8Uu
TPuVtELzSKp0fUMA+0QINSgl7Y3cjGV1DlbTFdc3ocqUxHdrCktAfG77e2VqiIoL
65L5sXtENr1tiy0PQNjuhs4WztHjfSjt3LEbsYQtr0huG7IDTLcZNAj6XFiK04JI
dZnhR2N/Eh6LQC6LgixzGCDeCtfjBU2EGkNP//5ES+ADrJvxRqpcxu2/qUd2pQIO
d4C7zpCAVK67YfoIkZp0/0+2AO+eql8ZUlt4G4554fopAlO+VMRwiwSHdlyQQVVR
Kuia1A5Buj1piwAV3ygQlt/AUhEpJaAbq4MzzcuKPBzoLpR236LD1uSWU3hHhAWI
Id9yQRG5wXWtXsMa+YGAZ6hGWAHtEg2u1IYkDzcKCfxIbuyYP9CWYcIorxw3V+F9
+KqVOu7hxNLOALRSglaJbquwXhs5REeE2elags+GKToGBjcv+PSifRPmGqY4Cpp2
3ptyQ8pf6fx38yoypS4Uz5ugMZW1xW4a3kGYWQDs9zz2pO7N+JhIBercOJW3eTJA
5ZieKesqzARynF/FDRcvf9XsLll/t6xASEcfgINguJd7L4E0ga+kgScFAa5RV9xk
Yhla7QEtPGe2RRoLmPVxFTGY85euvQonxdnkdNbh5ZcmNtmSJHSEVNab7vRcu/2W
dWxjkgeiCx5vcemvfpjMwD6Tpz2d1a/qZM4N641t8/z5R3nJv0+H1L4UsQcuZkW8
6xfVVQGMA+1urQr1kWkAp1tA/bMVmANbOyszTCf5dl9+1XapyIuwPoMH9maVDVCf
VqHEQHjyGxdM7DFLdfEwGnScaUC8LMcfVpsM/ufLmQebkhjH7b91UwQZydfd2Cda
+WbD9H/n29ryP7Y/phq8mRpExUtaR46RkMXDzbgAutuplpQK7YRo/e4T9HNuhB/a
PZpRxzMxAL0MZAM10fTMy5vEBkRsNb+B4nueeWS9+o7CRePCiSt/zcKRi044zqao
X2G/2CeVHNBuWPeqkivGqfRJqQ6MkRUi3VWwI8CNaJEO1jzaf39B6uNXhhRPY7aQ
9flZl9D9On7ZkE5oLSyTedc+AXsruhB7Lx3PsOJBeyhQnDYfvCQkQ66WmZ5LXs+B
BIjQ74UQ5euiAPj6R2bJImLSQ2a1A8j2uRP7L6okc7Qwr8zKxTWxpBRg3GgSMIy2
vbOWQdyIRn6Xu3rql1Kj1rEe6vdIHIp7Lu3d9NFZWiRVc2ihEs1RGdW6hbw7e3CH
RwcHlz0A/xQ5+t2VrJ/wHAuOWh6MSk6Oz8gTkpJhTbcrOAW/24gIUUAdXUlmhCRO
0Ih5GVYn3arwHWA5ttHoCYVU4BYF08BMdhbzmYVy+IDqecGCPcZnZ+4O/akHqMRC
JecsGeEMLofzSVVFW/oFclH7BASZX1uLIANZQ9jkc3RkgieN9F6PPYqNWXNX0+g1
J6BGpWdBvUv6LhroeGZ9og3rBBSR6bt5pBlmkc9fWp0ELzbSuE33YB13Fv8twfMk
erMAN0dGxRaRdLN5oYW7v/Je6KEVUDtZL6TS0syn32Q5CzPTzMh7KVVKdjorW8pL
IxhIQG4huQzhdu6wBU4hDndaY8+Xs+oi0+UAjQXRuDz8gexuCaiXUa9pNr7e9F5M
GI1wrJkDLZAb0untapVByGL9A9788fX2l2V7RjxN638TUQg4Y22cRiOg+uaO6M7e
BUys/poO23ha2LSvpfvon3o1qhJXRn2euMWkVyXhl5k76pInHrh4NAxantoPeTC+
AFogIP+QzfpUsWdE0H00LGoWdhK/z5/DFteIXeVK9npXAZdl7tk15PG8JG1UN0jp
TYS4LPsQC4MPXPBnkv3JmjN3bYjpnCQRw8L/5GfN2VJ4zvc8ESu2IMbq9vFyHE87
PNd9VUthdx3I72xsiXsQ9rVhCb2re4reG5KAuShSuCRjshLSY4nZY5Ug9jIbcTEz
LLwMwNQUMQYo1SO47jCK6weCM8pkbaLMhvQgNYWfF2g=
`pragma protect end_protected
