// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:54 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ZVF+2DvPxACinjkJnGG7I4sxHefm09poVq+EAJ9s/d7iyaMmxoejGy1SZJz+G1QK
/MqmBLc0l666Bg/aFJ85nVZvcvblEpjfkevSVnHCHgPPcd9VWS2EpTVRqou8CnVQ
dNUyYqBpskzDdb0ZjNhMrp2j5r/Cg+D+It/S1b0mOls=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 24192)
fehLYQcLbquXQUF3rfnG/NNRr9l93J2hNhoyyEpYadnz1NHDmY99lRoJBrttI4go
ZMvGS/3KIa3aIkcenhRwlplw5gPzTjKmRETHBvTn8MPTBoUIwFb+aUNddtogcPsh
DvZ2YrfBEU3ZXpTFKyXaoCB70+KueQ7nLcjuvcsmZPjWx4IyKISBQVfR3Dp2Y2WX
VQXPvb2JIfRRf7BGZpIIFjB6/wZkm5kKWyZMZ6xZ+tA+LOGJbLuC0IxLIXA+1efM
WcS/+P/5oX16sZF87goYghuTNNwil0FGOCKWJrWDMYXEsec/ph4YHg4dGKPgzCnH
GB/EwUZ2pBHMR9GtGujwpTh+9f6TS80pQAPOrdI/8WHqXeAI/EpPV/NvZH22INVk
0x9ARIfNP+lU3/ZHRdOYW0WlIT+unLAPYn27JkdiseeuAF6R7aK15rksGK88CFB5
GbZTIbdUlb4YRziYUhjStzF3bkhjpJT+dSE3FbseqAR1mdXIvBFbmpzmaiBgPsXN
MFsCjXPiAGzsUd3JeeTMM8Wza66qeLtK56de2z4P22wYJvjxSVjm8MiM5guZ0epJ
0HGgfpNbCdbQ1+NxhcVqx+pnTiQnFS8QHuFn6rC8UeSm1rFdKOhCvNN7esIiwbTf
oijH18fxn2qslaQOoWqrDfwD0FVJe97WQsxxOw8uEXJ6cK/qC/ZwVndO88pXyUL9
dizHMdK2uqFniOUPjeBaZPMrXv+sve85usSvTU0yeUqAPBnWaa+WUdBO7Qyyv2H0
qh8nJ9OHf8TY60/+xzJm2nwFa95LGuNJGWAkZ9/rB9hVltkSIeSFuTduOJisD+mF
Bl+rx6S1ZMo2OxejGqoYFvPT1BFgtufn/zEFw9/0ojxy2UYeXF1f1KK2qnuK5Vt7
bm292Gu3gC1X5PHUlfGby6I0zjGhRcJqVUmQBDbtd4U2whUhf/4HGpgbL5XlY4nk
Gsk+B3Ffm9WxeOjYXadE0jA/N9zNY/6fvx8DWEc9JaTQHD7bED0aj2tlTDTXgiHL
guAlINVWy3jbdAW2U63lRk2RW77yaRvM6y41LFbLxsF05xPt8tmPodC+X4pl2yUB
TPkYVktrrTVRtPyuocLq4uJ3b2A29m0GfFxda5nanjb+puHLp2yBhOrJBjLOtC/m
kAd168ngdLnA1y9IUsfooIexACloX+V1HfHdVvanlGXQGzdCDgx4QbA8OelnZd3S
Uhp1WVGzvGlrxIhVkjqdW5wAg/kLUE6II0wltD+5cx2ZllYYLtGolm7tuiuwWeHE
5zEi/s5+6u5OhZv2+6h8kQ2/S7bJcK5J+sL7CcWzR+y7RvYmyHJjvpYq7ZKnzy6R
QfCMWftEcq84iUsZo3xCqEneLDmZnF7jjyQKrpIhX8lliPOGKmvKfCuiFXZPzvvX
D2S4I8PJB3avRuuTyytR7bS/hA1k/GSjPUfPkdylS3DzB/DP3KT2CXfP0M8Lmp0d
2WL5r8TVNRz8hv4KEmhwz4jiz50u9/1sE2GoZ0IVvCO8cvWqPpjheyjzYt7nh5QT
O4WXsHCqlguEdCMdYY8hbfpwcakmzJJO5XJRb1Uzl+2UsRJphg76lCbwyzF7WxX0
lznw3hYEhxKHQO5FnxxZR44hd9rczCBqKXXx1HoQ7XcsZ1yFJdvbtX9Rnsh7JxdI
yCsM7fzjFdxskLZBmi2KBFTPeDFy9E1IP9e2b3qoXaVwDZfANDbmdj/rz8SGeZr7
3/P9X5Z8e/M80ekwL2kKY7Sp2892Uh352rLcid9sF56w3iYSjKHUmMxebP3D3tof
2pDZcUTbw7ghnC40okCZvLD/0v/KJoccfm+le76ZZoCFs8uOsZbuc6gdjrUhhdAA
I8fbVqeAq6xWVs4NEdz4hLAaQFBAGuD+d+LGVHHSbFVENy1RcyWxJE0Tk9aTahpi
0hx0yi0CQ+OaLNRzT1/Jvpk0DBxGZ0PobaCPGUEoS5ZI4P9hxL4Ugj7xJvoPq1YN
TF22GUN5PMOhJILTiZ98zGDBVXb28ElC9ObV69YsAAml2s9Fp3g0mA65PtJ47kXS
mSX+zqHcCwclM2ZNMLuuQlpKH85hs0GCZBpBgvOhA58bMsk5XKgr2DVEPQJQcvNl
IDyuH9uIeteL8zIJFEyNQVWYTT3pVm2EapE2niZPxhztUYM0Z6GMuWfL9La+FGUz
kyG2JisSrGM00tTcWPLmHMvM/tuYOlNckqWfFmqkhEtv5TPaSlYGe05zQCeSAwk4
Wuypo19QpXejnh299XnCZTpLqZt41CsKeeUWcV4KTeJ2VinmfpH4ACEkO2i/BMog
n7nTJHyKlvo4hDpRHS/JF9kk4jQF4bKvuNi/7Nrnt9LZaxEaleVj/7JaeJGljASG
EP/gYcGbJeiTw180838cZUToFojGz2j4HEJE3l/hYm6cBq26U8qn7BUrL5wtWgTR
l6YENsew7U3kmw66jGjDQnG8ZCY95WzAT2h/uBQrSYLK1QskxWSKUSYUjWGvz3ae
V9TCRn69bFEIYHIYv3Sd+QK4FXKOwJz2aKBCBVJz0pdSejDkXo856JJXf+wPyRA8
0mm+uQXZX+vajcYWU+LFo0zIheSTtTmHGDAPeL66Uv5MPx3O1MGQNNflzdEjOb8O
ya+F/sy+VYxoneExy+73FeRSxqPHcPav8nQV6mfMWJdgInO9j0wqF2/rUxk8fidm
Iw03s9EQbwpxdF/5kzV2NMH4SJhKS+0aDMeovkObMpcSR5lB084RpHYWsZdb6Fp/
of3Muxmv29nosNMsT+JDzpPYpTsvVFX/BNkk3e7Z3EtsxeUcTijE6DTIkMDYZ5Kz
eDfwk3phMBuEb2V56G1ndTGNmfYe7Ai9Uk2Zv8qXLNSSKHP+0gCxFpzwk+K7rjfu
AJhjqyhjob/OGoYfeIERa4dJMBh0ciPGHywYjXVFpvCc6yO8eaGxOtkz+81RFECG
7bfhsN1lGLCZRbvdnC93sObn1gj3WxW6IbwWujVVskEqM+1YeKFXG/DcFrkEZUv8
dy6zloRsb4J8StOvtANkzSI62vfE3cedmpHD5gZwibNZXBo++3D669DxuDDoBnGF
9v3v8clMlIhP2NOPFaL7nO7/OO9n4MrUiV0PeLq1+PPOzMlCkypIFuorrhiklSVT
II8mGP+mdCygCO08XUrnPCvFq+LVhaAno/xCdgA6oBI9HqBqFdT5VBv+2Ho5LY+C
yDs9VJS+b2vH8LFq+dnvdGT3ngzwcOSy7m1LMvQ2DfxCeF38R4E548ad2HK+VDhI
8ToGiu5XlZeFTa1AEzVW406hDJoAcloZAJEqBxwkcecbsvz/qt2IRv6hJqynDiUc
RRW2oeeF+LMEImQ54CSxxi46PyU2NCgET0l3ZUn1XJ5ZsTOLFEA0WPTSlTLBsUQ9
noAXXUe+FIHyjXCR4mOnEN+og8MSk80esGM86hsoHhscvRfS81IByyHBYNUKbIg8
fvrM1xI80evS/0V6OwXRB15Et8Uatp5GkGt5/RfpPkxLaFl8oExcStbCHuBw2nFP
M9ADUSSAd9g/oXu/1UrQ/HsrGFUiXU1+ipRIsDgk+gbkuksdbmmKO1as1LET/RXy
KfYR/tazJdRVVCVEk1Y1TlxeHxHytFZ02mvphfGIGwSzmgIpvpM4Macy0r2MyiYH
7CbHzpluWkd8NHOYEFNgOue5gNAq3DTJwRQscL8Kw01DQvSc23YOGa+Jq9dZ4acB
l92sOmlq26kv2M5HY7JiOAlt5QGTeaf7UmeCGjCTaJeliO+SKGK3ys5VRwRyk/Mc
puwJHJaI2pFGV1Sbn6Tkgum8DbiMoJLO9V1DXJ4J7IedUSOyJ8CV1T2rPwrd9D4K
LU9zzKS7QqZ4WB7ck0KtL+ig60bi/WUXxwmk94+XPF3wWtDobSfgMTgSekLnVjLg
5z52W6yjn3oD8UBmIFmTgKJUEujVCofDsZttVhXtYA+YkwNMtmLExon+m/DXeCHl
dwUIG1HJ9rrIJS+jMo9f008CJYPXh4rHzg5anvrhHXij9XOmXIpJ5h2bZn0p4Wec
/TXOnC06+lbXwHihUCoBZ1rMW7S4g7YaDdLRPQs6qVh3fsiwGGA15yX3vxW8QjkL
aRyuzv6Q8BhGLBVVtvyPfghvwKqYS1646HH0c7fmX0Ubwq8eP+F7SQ46pO0TEqHC
W+/tNGKJNEh+BWwK1nIBYfBurmHGi4qd25jHBRql5H2dkD8Peova3PcsQE/m0Ua8
fD8s1xOSd9opRUJAp7QkzTExzpYD0LJ6BKZcTU/iPzTeWLSV/Z0R5905SJtESzPv
Z88A+57yyocEdL79i6FMaNNE9LQSQ13EucYzyQv2iJJUR3wuxtjC2cykmtGzHTNb
8RXeH48iY/IArPIJQTJjR77dY55tShkhp0OJhsLo7FBK95ckHKcHzZ0amIhmDDif
YP416uW/dUjvl+BrWoh3S4wFaqXVR6IUw3aS0uSfhrEqBFz/5tSN50P/l76H4dal
3UNUfIajqXaO+ch5zJdfO7I7dnts4Spf6YGFB3oV3Ah8C35Et+dMi5aX6Z08p0fo
xN+wzQk5bjWpstSEExURUKbPBV5s3NK4aOoD0bRTDs5XeycG1jPajgjaiHq377BS
IqFfeRfK8OO1sOQi3FybvwZlvu3NyX8ortnBeODyh/3xEYHsGiHIx+ceWpM5Og+4
3XOYRHrj51lTgGYVBLTkjrcLGDF5pBUG1TQOrPOlYSS3zHUrMRkcb+czLsmtwxSx
JTsjA2dNdE3oG5qMKjovRVQz3SMrdeXNGf8p5nbsucC12G4uy/GzWSi1YA6/h6L1
fB23YqhKhsjAJ6xLhXQL99mZqmztHVh/AzkYkHg7krdDEUyZK/MmC2WtSkm10Sh0
5d2pQgeBnNSxFnNpaXqqkTwEW9QER0lq3tQtHaRsiM2vVdXHotcf6fV7r4tQNvSW
BLGI9KhPKA19+t8C/vxzBZ3se9JCR6+Df5d+RYwLa8lp4KPC+AmM1gbP23V+kLug
pQI/D1pTOXs1uf+BwPRRHz4gih0iHNXT/Bo7SkVp5h6tfOceP13HLwGaiIhPHtCM
hulPl/36HgO1y7u88EvPoW/74Z9w8HgXo3gG9IP+q7EFu8j3QFXwOE/uO+DcnGs3
BnkPnuz2hS5JTze78ltHxjyB5zAKufP7+FUHLZQ2il1wFWZKI7/3hylp4Y4FF8dV
ZtPJVMDmz4HXtOLB1hWWHLuZ53Pl8UasASeR/afDp7Jo6ZWZZHqoVN3E322p3ata
tq+2PTHw3kE8IKt5dScVi50RfO/Eo88+IGZO+OGfiY2rLwEPyrPMxXt4XxWcgvWS
ob2TA4M3t88/4yH2iHxPYkUcvnKBzR3hV7fJO39LYM7hZ0DfHBGu2S7nw24sTCem
L4+hhdNI2x3/wtQubKxq8B8yt093n9+lt0JhIJGfMG1quqWFPe03Ss0nPheXdEuo
Tar1fKqtOZQnfMuqtxOvXj8Jo6rarIihmXrHpWy2B7WNtUsZYXUKhZcaBeFqdlUf
TmPRKwzivDsTwB1JNE7h6Uv7XismF9P7ZKHtUpF4E/vOYLLStGeM8o+b/NH6s7pH
zsvtWUK4FK1RMBsr1OqQaIwiUdJP95Lehxm84hasqMP4yV3VuNOFsZjKumhN9cwx
6LO63yhLLT/00o88DqcHxydyjiuOQgCuyHX4MpWlbwqq/pRJmxpT5B3ye/xxi6kA
3PR1lQVeJn0i19Z9f+qgZg0MxkwBGoZkGCz7oXuntPfEfzaMi7O7cJjKBbdfXWv6
f6f+QTje9JZyUDAzE/m8latp6W80J5nm3SCvGnfFc/g0Vlsfy4l/WiXbLTf06/Jw
KV5xzjx0kNk7X9n/+AbrCmvuO8eK9arr9rOdtSsvzgkcP0OH/13CNHEtqQkI70Mu
pLHTGIr3XCw6620nFJK2C7pRMWJZq+o/o3AAGwSSA7+2RrMkIEZAl4L3wvIdkIrB
sd0b6KuuAY9Nit85AGlQGqv3sCWjLGSVIQJyuJPtRR2aSUJlCsCrEWgQcQYoNWnC
4+W38TSFHEzXYtWQiKsxpm407dN2cOmal5MBc+L4/xVGU8Q0nsNVn5pyGzgG36h8
g4NgFXzxK7Obse6poSe/CEh4X2v0f15WSfM5K/hGyx/i372plVKo2A0cBBLpW+CJ
L73XeLZWWME3vQctFtZYKZ0rfTq7c2fIr67/gKxVfCmo+aZu8NTMJg3KxVDCuUh0
qD9tUfv4CbLakF04YfhWnTQFyagfpuMtWMh+pW0jLzY7o6LUnO8RFVwp6rQhSOQA
2BcLvORyei3hi6HzKU4msN78WBb9ON/gSL7mM3bLfOcgteDnytT0XJHbqmQiKNjF
tOQwYS+LMaLAp3Z/g0L4OxYtlvNZB+msXvqttmSttAnPw4Ecvd5O52f5KKaDBBou
vb6oOSR3/IU1fkZ6sqbS9HARcSRcQMaLLkLOYfPGAxmvQjUreYOB8x2IUtcaMtLm
GKlbFvQekCMVQn6fcmhT4vPR61koYhqneVjqeazJx6AwNjemI/V76yM4tJwYHWQu
bFtcUZ7oVvwp5KpZtFaE4Ti6ofhTwk6yUdl2aasg8zianO30O6LxuD3oDHAvj7QK
2wwzSV34BVDZKZXRfJK1SQN3HOoTTCX+P6KKcNmKQqsYxADdjYNS57Fi8uc2shry
zZDj/XsXNm9zfd+9NNpHAYz1PPQxFP4NiSMGFRVNL/sH0o4cIoCCK1mtRzIkBYSY
qePBG9Xd2ibaVpF6Q9cESuy71DeXuPB2M4AMTO4NVPwQzOMXRvKH/ePhHNYfXgYP
We36IFFRoahXTksp92rm7X2nMVJlKq8Fuv73a6P3pN5fx3T9sDlE4fWCIUCM+vZb
V9ey09QilDZ6baezgoWjwL0DRG/kGrD8t6JzqbizT4KZrtqq4pOpbz0F/diHwi2r
5rU1R9X1o27kIcX5/RnSKXxXPr/7wuTAZfO74GMmOxtmwHE5htZDotMhg2xCMxXL
BzzGSzb/uIQxiQ0ZoA3RN/6pPzXn4tZ77rCq1J2HmeawZvswdn2yQuT6ZFSDVesP
yc1MNd2n0L3dRgFy/pnQmLiFMXTBNlc+0xYstCy9YBjldqoAM6QJDHkEJX3ML9OD
2u4OUMtj821d6VCbTLIp5UUWTPy8CvJ6HhOHMo5WXsQw+NsSOo4pcK8VRpuUVRs2
1+dDFlwCoyFVA9poZQUYR90pYM4lxpNABRJLWlbkH/0i+fyxW5vMrAyDrcnuXl7H
5AIDgKMOM7L5xfzGzR/R/qbvG3FfRGHxY/9IwQdI5T4Dfs8MOuyz7aT3i2lSQ7sk
otY/CkKENzjYI5W/s4pRcLtEYeq3eDcAtp4fVApcdQp3tTq4KkLYpXyCMcehhWDP
3PW4LTb9e9BfqFX6ZAhxvjQNbe8kv57yz5t8gE3q160fAfkmSMgcpMCezwtFSvhu
6ELKTyi4g+WbXEZLJh4bVSjVMc6yQO9zFJKN4UY2Uj4qnB7/dvlmv9Ketj6kPWQb
pzmsFhMFAYceJrEKeMG1X0QA9l6zW5TDI08f9nshJ2qL8SHHI/S25EYvOh8VNeXm
7YRo79LObukFIfh9yH9BcFSogBOyfHA+/6MlBNVxlnx+udz1kMjkiw4aYa91nTen
kA2iXiq5PhRhLg0abduDcUr8VE9jJTT1NJIqTtsx+pcohxjwi9Juzuo074q3GpoZ
BL1QRvmTT9YUlJFewj2gIa1JrKyw4m0vIlUwVMPCHFZ3uGYYUBEnIdp3SDsK30Yo
mbHkXCf9GJYriPZqhK//P1tfTPNQ9C3i/6pdnt4gMItEwzJnhax1/l98WhkhNKiN
DlsAAFN7WVoEBaIKvWRmGV9c5XO7HQ6WPHGA5WgWGjyQrxzxPaLQPt8Dn/9fifzC
J615WW9CHlGuoh4CbLRV+HsV588UUePgdqBY0aLd9j9kvzzJ2uwN5c3lzzaA7I+3
fWGKUvTBqfbb3osNX8HFX5v5f7VYpULjHkGw0K9Xnf513CHs9ikroLKUibwcFgat
n2F6nIWXpTQgHnPy+/pFmxEktrhiEqe/KkSdQfbx5hAGHT0bEVwZ2CxMGUv/ZyC4
URYVycZbPxmex5m1aom97tb1tdAbEw+H2zhATufCMoamuHMQVrwnfLxViM0mtjVI
4g0YmSLRcbqHFMfgm63QIZrhrSjyhhu5UETGggGuTxCNFp33n6faGa742wO/7oFp
01FKEIG3OYZypsg9NRKzAnk3l6uWp4h66v5pt+p0w81JRsue2kloCsHvAuCmy+Ns
xvhJ5yKNyd6m0m0W4M2CGY5dZAJs9M3NW8R6rJbOxMrtA4oDDMW3mPVg+dE7mWPv
b6dxc4L9irCxloY2qfGKlVhQJJX4hI8tW73cwpSOMRgHEZdmrj4bd/bwHxjRWDkg
Njpk41/SQLHP0yc6woPvWoLte+ihAXlpXHm5XmZWRM4mtjagDrPAU3IUNr4q9Kdq
kFxkks9v5i2AA2kfCnT2kUi9uyw0lLK4ShBQt8MmlHCUhZoS/CWNTaYPuBHJdnzo
/yIjIZYWopAm0/Y6pE4q+aSWYmBu59ZB0MuoP1dvHiUbLh2p9tXJt66kc+CfZJ0e
LnXlXcD1tMueVakIZhoyqMV0ztLe+BwBncoJLyIIwZx5GiYlgAFyhJL0Vqx/x28B
aLtIlKKBSD2/L38Q/dhyTQ5VoHlGufi4Ftv4cX3YiPJg3GituMEvY+Ak02/QIK/Q
WubWSzCtljU8WsEPxy0WFaATJD56/BzT1i5Ji3OStXqkLlXYTeQYY0+h2BfkQBP3
1kDVdoiyqVYRqIzm1qIMNk6ydscS386yg4+BtkQHlvnb4KG8ulfWCfWizCXlBGpf
524g2RiWjxiMdYsE6tPjUOIpBni+cNRSM2n/49aSKNKNHiZrN9guIzrUaHv2NVIK
1pehvvKxqjWM4KFQCYwi5Zz5WGXqor88323S4JnfOoHSfzbq+GXDpLcY2ZginktV
5DfsgJP9FAE60y8Xwy+HfyqHU9XgjlmhVzAgNmhJgfZ83/RA67LoAHVgafDqANdO
0Jt8ehEAUM5MzsEfYj1FkM7qSS9/OThZNbPRswG7j0HaPi4LcEDuEC58PzBelp10
2LkOrHy/5CuLJvRFKnP5kR5FzH7IyQK4ATylRzj/5QIF9uUVMMWTsuTVsP9KgR3A
jsN1voIZiDnYFMOsHeqq8NkDjTS7QlafXdEmUp2JMZ4KnNeftZlbboP1uhIIK+d+
x0t7GIXXRev/r6RlqBUnB5gNm4IolaYTRghZhNuoEhaWkT3eOJVPtOFRdS9OrK6y
L3GbaW3oT9C4wgnr08Gzr0thtj4hcOzuoVHO3BS937S92LfmJZSxGnolj3TzsjFi
BKVg/bAJXM3kUG0Li1M9dAU9PMZUvdAs4bGlp2ERrItqvIYHrIp/qmWCtCHlJO9+
V1xxHMPOawJFMhZ1+QJOtPTMrXDUUUJMu+ti1rMU9jbqYqwF7VwTxyk3yomN7vm1
9yW0sbxHsGoVu050X5U+MBOUZ5OljVbcO7WffnY73sbPUomqATjpWQsZmo/3fMip
iXsGA+kpXgtQrKvmNA36w46GvMhlhZlYCapE8riA6BHKzv0rTBtVNtVpcly9aDpu
jAjJl7STQLWB0YCcKQIIFnmu6vdZdgogZot78PRKUnzgt88QChZAwj6TLyP6l50n
RjAmw1Z3Ts3Axt52RUgNWo82K189/mPvchopG53wC3u4b6KEKSQQJbwS2PovofVl
v/EOpPlDm5gSdxdJqf3sDCA9Ym9eWMF9Wei1T8fO4TKcLdsjafouEOXPjaEwZ6Bt
XaX1bkLT7YN3TxG2qxGpM4N0z58JkoIZtCS1TPKFr8GZaPFHOcJExZtp/bIKJFZN
hc4GrtgJy4cRydbFpYANBaQ33rEEy03Dz/VGKEzLd0KPxIv1g/5eJE2VD3/tkD0d
sPN5DQaLUASHC7aFVIQlhLDV1eSF7Rq9mH96WxIBnaxb5rop4paE5H9a9z9JpASG
BPHgE5/xJ814Mu38+P1vkPTnTWXn0qBjNDNYukeH86taOUyD4FMh1ObhYFvzSGXQ
ZxuDH9L2hidZwG9xxxd9j2Ugt1Q3pz4nZqyeSduVn9X6/HabfVNk3fsgi16ujqpb
xYBxQNaWBZimZwMsV5urFaIp28ShfxUsl4TO0yAbVg47TOtZiNf8Ygz54xurvK0U
JbGfnioZENOfwZBKbbYxISJkojDi+7Ux5Kuvd1X9R6CXELp7qhT9hFE9SxrLRiYU
DWdj5YqFADD5QXIEubEUNY6Fh1hYlN4mhTbmGZm0tJHq5OnK/974RjgX67XbIhCR
pEuEsZWFJ2NW9sObWp1xpSs/a4et55HHjW+Xt+oNF+VWEZweJ+r8ooL71aTwlUYW
v2hyskuUNWV2TErKV3Aaqn1zhvjPjnxVoM0X2hQGIFWQd4Klhq4r9q5CNYZWoSN6
h/H2+TQi1CQDoaby0VDFVjCgG6DSWZRNTpuSgZbZEWC7WlJS/d5pAn1ramgtQABC
i5+AAoBNsfGOObDmvKa1nJ7pVltAOflHftYWjHWMwqYJvNfAFgmGVRDAbms7mvyA
rcAncHQzvpnxRx9iKQY7F6R5W1SpwnzkzD8a4325/EkreHncATruwJFC0ZvXWddf
qM4uCDWmljN61Q+4nJamkzEXpf276i6PTerHrQznF2nHkmOJ7/SH1mxKoX6zhlH/
6BKCVAODmN43ZjV/cKEuKf8b0f3qKfhMVT30uwYGA7N20PBhrfi7x/sMZFU4LpVy
yke0u4xpg2xEjG/w8IEBROWT/pyrYZLqGswfdqX/W62GP6LUVpxkX9VEyE5EJn/z
FEOS8gz13x9c9GpkqQ7E4v0oatD5CfWktpUc/q04U98zqXI1w/XLPAVVOH94b3t5
BzEKVduqtSe3RNtBALivrDEVZ0igFdjdflc1+OKtdX45CxwX5UsH10GsBpRy1Pqs
0amq55nszk3qPhPDaqxIKlPcOZsUvLyqbuiqD4wSMOPYp2bsKL6zUGipBWOkZ74S
jUS8IoRZmqNfCEdwtaM1fNp8hhF+yLFFE/3YWSYRFUeitGvuh5GYiyb8L/pvKmlc
aO2IrRsNHJYlGD54QmWMfBYZXzM6shhIb5ac4mmrN2mqXwnkNch8BwAR3SLl77uz
leqB0wlOD47wEsPBzf/iIJMmnaxOrHxNVzgeftyI5L2j4SxaPk0hlMvpQ39pXqRW
1JoERb9JJGqVbn7x75fLa514omxZVkH1BJzl5sP8S/T90fUVUUwHVoukcmj6vHby
o3FDR2VWr+faqNZ5lsjc0WurkQM7kT/QigrrVMwMJbwNZNWJEwfnEqe5MqNZLjHc
aoy+eJyT5n/qfq1FmofAKbBaBDGf8Wzz8d1r7zSuOlAmpGg2UW11JDwNGXAPX0ki
z5mmm2T8BI8i+F849DeD1kJb1Q98wUzovNYav2cFwhhq936aJfOreTfuWZGIc1LG
VvGkc914UmWICJyUkBCrwwamPORyVn5P5Tht+QN78bWncYAnUfZafIqMPQI7Rdr0
f/jPKReQsZUjacZvpckEMcrqC74hEemld2HBKLzOQie9z3kpwitWG55BWemf8df6
pY27DCw/bRiSHe44GP3STUt98a8b042DHrzMqQ1hPeHz4G/JS42xoxp5SNYKR9jW
eSFrLp3iKG+dUd9kV6+Vmx9hFnMzh1v7ZBdqqFAwvzvOrvI/nPzhW7xEjYF6Bk6u
ex5Tlq0W0+MVMwWOPf+ici7F6amfDA1Q7R2kM9FF2QBCIJrl1mmmDdNjpdO/vNER
2g7zxXSYz8T5i5tpq+AhafuyGfQa4UxRT2RHAO+fwNsbVMoqsWnfE1O3XViIHoBy
a9VEUMjGlrLL6wEc63COnoSsnfQHvvlFiJ8BMPhnPX90WrpSPLvgFDMnKt/T0DL9
NQ09t7LubHyGOQABhISUKx64rSgw7/evyPVyY64fgeqGdKDeow2js88oMls5Ex9F
jQQ1W5XhaRO5bCYKQlzxZj2BuevI4zXY9CG5YK228O9GPj4Rrd682LFvcMAuB01a
E+P378OMnY3vQ0862XRAu1DajHNVgj2NHdrbQMjEGfUpo077JdtVvk/DYasJ77s6
waT+Gkn7pxCtGEcshvxg7rlyoCvrHKApkKUtRWORg8tG8zSs2FK0nLqwz5q1eem7
v/t8o2Svqnyzk0ZFHLa6zBhKVKHfD84mGfA3LzPTNaFtv5xNDZyZXC+HvfZ8LCzu
7eKlsg1l8+kWZAwkqLOGGpL3DkQ4Mwuza+JQwr2z6IcKfsZN0UutaH22vijAu0Ml
rPS292n0OuP3Z44Hkz+5jvC4eDCZ/tJPXQMe9aKNgxFwXN6YUi88S/zWiF82LMXY
gOETYF1C3asz8pfc7pfzBYm4jsLCvJRUaLceU7mcYAll3MHkYoQ6h4aQ+ffL29+a
Ktu8XoiRWidDglQA3sYJ1/DOkte4XnUsp9L0JrjyCs9yx9LhkwDcmu+8zMBz7Ej0
sSxYf5ZQZEF6pzHxyAJI86uXUnYkH9Au+1/CMnqMGBqUhHoFUi2pUcAIm1s9Ddta
9NULKcdYOw3Iru93bH0S2TwYBeq1nvUfxnqSW9Ww7Q44447GMpcAPd8nwBteMhjN
J+GkTNLo3rMP2tqfo99yFHl0aTFfvJp0esckmnYxA5BcAhlK00rvPVQKyQG+nFze
d3jDnOQzbPRIWAsfLI3ferbn2Nflq6pi45egMAifOB+Ezfpy0LXWHWSse4+SBfc7
mvrxlN6M6GB/tr4jlnG+N4npqzJo3kxWRkcfQ0uPgqEMRyo8wxtph2lOb20qRBj3
m8Icx8NcjM7ZlOGoYnA61619K2qPTjJmfKec4XmwU2hPgJiqmSpJ+y8XWyapfQOj
RtYrKDNwNvD0EsC3KLxF7OnCq5c7/0EeuoV9WpHL8iT8p+tJ+TBct2o2PxXRkckS
CnvSatBm9zmejECQtPbsla9t/RdMBWJQFJYwz4S9geWudnGS2y2i9O8ORt7ejjHy
xL5M6Nfikd4qVb9ax95oXY1ZCmicCr/WYHqgkhszMEvaGox/OS9rl6jsLMt/xSYw
sI5lJ3aOLOyyln/01Z1fgHZ4z78X6cfoesg1uHAffKr4l5+rte0hOfMXatshzl/y
IUTcb3ojgDjzr/VfNA6Gt1po7tywqeTPa/Z9AgFsfu79AYegwflIWrxE4QJRAwxM
QNErq6mK3ne0AduSr61rUBY8cy3iy6rVncQood08JDFBbA+zF4MYueS8LJq7fmyD
dWz8ZAcoos531ZHpMgbBKLNPEqdGQPMMYsQyTXydwIfnPL9P/09knBPJvfX5K4gc
RXy/6HtbygfnV53eD8HIZiL256exO7I+i4tZh1IdDD/0w55wEn65WoPv2KC0kbm0
AF1bIhq5PF2B6CSyi8bvaPDsS/BCFHHShPRuIF/H4eqHMZ/MzJI7hQKr7ZbVALU7
IRbci5Fi9JSaVpNx2rpKbvjVfmWwbXIYx67zJMwePp+l6uXMC/aiHlrpLl92SXLv
4EvMHcJQG5kuoaT30P9Nul0iIOekIy0+4nZYw9EDd65QvQg2XamOYuU+v9XZDPwP
oKtImpGADwXG8Lg7jKUExZOgOpvmkz71LAPExLLMb9ywqz7xkJi4cUG2LKR72Mmq
dE5vE4lj3/rhd7vqBPNveq4IYtAdrR/VHqMauZsdDJfCO17J0OoUcRRPwvotXRIq
f6bi8ZSz/lexEfY4Q+hRZpmJ6uvBEnVkyVhPei/l6r6ZbKjOv125n4JCRRledfUB
9iifQyN10MkyLq4kw5QhiwnlpfHGmBws54aC4iebhKY63FUBu8N+Xb+nEkD9L1H4
4FQhoP/KwrWD/HRUV8rSR8qTHr4tjpIY4Te3taoWuajSDcq84qnAMOM1GhQhBDCJ
9UklYRQyQzO2hVLHzumx5TYKJNsZ2sH8FazW4X3Eau0OVMkC2pKJuxl0JDNEveyW
rPC686FI/cyNjOy/JNliLi7wXIHm2CM6kRXuTu85YEGJSH03Buam8Qq8fo7oH9Vm
Sd1QxyrJi7lKHwOOQkC4hs5DFlcMX7iHPjZAoUi+U8zmApv2Mr576vk+LQ6tHgp4
8U0mPTJlvUGQ/IOKv+KhGXgC+yjYlJB7f8rootD/3+JcvAp5uA5JcOV6Ww/2+QsH
pvO9UpPifKBpKHV0DAgVU5zMZ/Qz/cjfiK4FCXzogtzzHhcXufHHdQ8IESSMnDUq
nfIvO9az7N5z0431JDtRZSFSlYzg3q1u+jeQNhgnb3Jh8ies0KT9aCDLNOhBXYyM
t3Uo9nCGd0duLjnEHNTL2W9XgZ06uSjWO2HTVvXTk93ydkmzgMYzg9jjELq97gJp
JkMdY4D5GJ532YPxz8nJB9lt2sx0Ouyaniq7HSbXCONJyzKDM+3LHBUaOg7B37ym
6VdwnCPFAsWt98i25brXHh5r2PmmpX7NvEPA30rhl41CzbUfA/z9FlCsudH63OPW
nvxbb0zr/45JfrSoX+s4EX95OABvNXqyWPxZ/Z/KWg53XWP1anFFhzCDeeilnmab
pb9RyqkegKKIr1DbJP60W6UrQt2Vh64fD2YOI/5J/91zZaHUmpFHEcmfla9hHNzw
uxzF1Oiztyyt/rRll38vjDTrgmqQW3XhFNtu2ET3SKMWFck2Ls2Z98dYHTKytvx0
z8zv3ik9qcvLGjshwYSZNdelW2ykfzaYWg8HCb0MoGk9Qcb3T2nrUNNiuVJH9Bx9
i0f+6p9WRbbjZthkvcESUmMs7tLp/BDPMNtwkLtgow1X48yJjF9jCh187XhjZmAd
VzhxbzkGYYm6rrUxx5CWYb9PzEHO5ADJt9iQ2VQPTupT3ZbXhFkxvindBIUIzBxy
OGwAp6vnr+OZDpfw+a1enfobyN3LyoD3GITiTqAYrM9pzQTJxQmSQRyOYHI8G7kS
1uybZOFPj0Bye43jjkDfrutUw2nr3kxqkG4MlMPp0QcoGaRuhiDe7uYCA7xHUJm7
XATuppd0VbRsKED37tgTtmRB7oGdjagpch5S+afKlPGssDvgTMsF7n68QjLor5X5
YHjTOTCeloY5gyKA6dHTR6sYQQt+wTHcK1N3SV8P5veWnBMZPPNU6CbN6n68ttX6
+OH/zsdiPjOKsMnBdqzhn/lDaZD0C6UhNPIaMtoPnSsnUV0+R/Zaks081OWZhxGk
QEaenWwft4d8lcyTzCdqUDbIkZ84TWei7ZDPr6V0lsJJj0OL3nkb3ltGwqN9UOFl
YWM6AE2rPZRXvx3+wYDANd5qpnqWq/aE77lEUBoAWBXgSIRC8ipPZIb/4s9r2Gz6
CLEpeXDPffB30a8JskA9x4ZRDbC9KGhtTI5Xbp4Pa7OTnXfdEjbkGr6KqeNyXs2b
co1XZQGhekP00StF0PWtH5SpakwPFJ/9HgOm4XbMhAiRk+NT0/X+pSN5aW9j8L5K
EG72qHnZ1yWbe4MMgaMYnUXB6rQw8VmEeeFbyrDFPCHv/Q6+d2bNZ5Ax0H2CPIv2
6OgRrTXPyZvtpXosYUDLHW+dSJotGeTUdMGNdge5nEBSSIHLn/KCwI1OFOj36wjf
5GYK/XHZnC9gecSqeI6gO3o/jEpFCp55UZncdseyg2KK5Zc/nYQvrkRbyzkeF8QU
eQUeuyYRe2cID8yr37eU38VfP3ID19snxqJskOqPBE6CjRomk/yFKJ7ElY/iIVaJ
pTjawhjnWnpJDLEb1ZQHvEWSScKO07/tZYVVQrOwRRX6zbPTl57WjRfpN9blkpj1
G6YxUydKcPPBdhu4PRW4nI3ltgMx6POuxECARaq9p1wifZV/7FTheeDBpyOpt7Qo
fIgF4zLVzhFig2No0WYgiSjGlEK5wASuYQ/auyvuZiyQq5jZrvl7tWf59Wi8GqGC
LRkLRMfZXsu9OYLr4iwDVA82q9Ap2waeKbJNE2v/hSRcaWQt4vqLII8G4f0rR5Xr
sd3SULarvNu+7YVhWOi8VLSD4jJNwemY4oDzVeLmM1GyseycMxJusjBDgIFqJNeq
8s9G8FXT9/Q/pPBX3NY+QApuy5mQp1mvg0khsgeW2QMJAY2uKKx0tahJmmJSD5+H
E7Vy1CtXNLR58etPjdEQtmeH1Ks5MOgI5h5UcxsG8X4YrGNItyHAsFJabngQEQaW
AsCNXn16nBhG5ORUb836y6bxkNSfrJFjwdcUK43Yz/irvi16mFVU15/rDVlAE55q
Md1FlnZDSLKv/SaRoFyPVrpdgNvlUQAbfgPp6HA4ezc02KDZ/Ztkg4SH0AGN3hk3
jPvxq0E2ctPb2GHN4HTzzTktegidWHpdf/ZGJsCuQl+0cpbsVMJp5RwjkDAcin44
8KGIGeJBIlvanvDdBMHqPZBG5hzQmnIkukYSejT0lqAVyOp0wm5Zb2GFsaQluhSQ
gQU8JBu+EcxFG+fg56L68Zm5Leo6CvkV9AnUozaYmXY/a3DCrlHpsUE0IQZDPRwL
YVKZ+PbPYt52t/2OzYLWb4gfoFCtBNhhhcQgObMafqGC2iNqyluHSG9aPbh+ZTie
LedKo280Z40ZPHUJXjkhJ81Ku8mYTSNGFCy7WMPmYbafR5OgzYPLHsLYJkV+rc6a
YOqqnIqXyYZyaTCFy5RbTes4JdWZICk4jntXo7tz3LURaWJIr60ULTuXXDEWYMy+
oNIf3qNfwHiTHbrBcbtTkoJXApbTHOYwj0FBCRqMq22/zQtiDrvXwBNISQ7VX3fb
OA7mxg+xrwt16eYH03De/YRkrgIX8patXasN0Etim13auXz6ykDg1ljsJNBBujhb
H96PUoYH9ybYpU+ivDKD2qJyLJe+vW72V/Kq/E67n5mzRj3YEyKcSl+4P6tcWbEz
ps3APlykYhqC9+Q4nvaOhVYyLyh1nP4DLXBYD5Gg+uVcHgX0Dj+kgYDEzrNcd5a/
tESPGFzL2z4PYQJronjcICEdCNbA60HOCKd9c1w6i1yzHklyHnyv7On9vqtKcpZt
iUWqsi8ob6jjDb7neyvGfiLeaeqOWw8ekRypaX6UwXW3T9YtJuIz3Biv9RcF2/rc
MCfNG4xp2L2aqPYk5ufAMwnv2rTwN3J2fr/0OLC2vJfAppoVqRwj7aHV9zDAVMef
6mGHas9Ip5oV5nLjFkn+oB0oIN7EAgVlSDyF9GauB+ruQ66dOU8/DAkcLAKdRcqI
RWWxS5yf1uf134yd92EEbG4vItiDQ20XWztSW9pbwJ3Kuzm5cCNvJhjdO0bN6n9Z
Kwj7knosoddvAf+oDpM6AHreazIOd/5Dz2A57+EAzEotNCVYLiJY1oaIVZovRc0I
ST558OKjJwFLHHFjnF3Ic+i/Y9j6V66IrArimqQotPc8V4lt4FPdWsVoVrXn5qxR
jmGlVpEfb7mZIuGFCQCcE1p5/26QCwmEV380Le/3CRDV+SX4uNoUo2XHCZE6c/eP
/DubBbcT6Ri17na6Pl/vMi4y2mkMm6XhmbuCG4DyD1T7TLc37bYWLwUy+MwAsg/L
RkmL0NMNV9Qg3qA4/eWd0W/VJAImybZksTeBs5l16ZAnwN9senWkBV/SCJLwHCAZ
x7daU1qsCE4BMaBkc/B14urq8p3E8VBqcI+3KtVfjWOXlo+Z4IfWRn/gdEk4OKtq
840RVjHGlHH3n2N8BPZzvXzkEWOR9aQN5Tz77GExxLOv9bI54zvGJlqSL1epm2kG
ktT/77o7FPZ0h6fMLJlhG0go5ZYC0jaisJtFBhIopgYcyY6VFcHPAkpmAxsBXd2a
gqTqhP/QPqaoAnYXa+N1wOQSCtZ6Xwgb4y82ImGbdsAYhvkejmQ9akahORK3rK6K
H/JpV9WnsboJiosyyR37pT8XFpYwolBArZPf7fyamdNQ6Dgk4z2lbmBHHAy0vVwC
L1PK2LfDGU+FM/d94HnY4sdsivMeXYOlb+wJjs/20Wlv+mWNnsLITIRLt3D5YLMA
bpNPzKOxis8dmiq9F2xZ1D9j4tfE1wFnJANBD+63PakJ2ll2paqtwHR/wdigUcrJ
AgYh/Sx6xQ9cnnEjpOHyvXk8K9B+q6I96c1hEQInBN+FTJqz+ogBJ3323P1JHPJt
DJsFl+GNEXUhJpeEyY1NslZ/sUYO4miyjMzxcT5YIOm4tFX/x0zGLqwrwSOOTKqe
9HrPTcKGTpWwrJ6uZTzMzf+y/yWCWgbz4nwWmQmDdDOo2P5IAzztZgDilj2dUEGb
FfmeAaGqzIl2fZSOumRl4YIJ/CuylmvdE1QKLhWfSgouHKZzp56zXSPrOA+0aIyA
0la+fa0HmcbWML92hSStVU3hIDbtlz3XPcyfubPHrFhY/5+Ba0ipQNSa/heehiiJ
1gpR9ptPiPi57s5ScHWDW887A+/W2jbAiqOOTaNwa/RYNJRRB3JQTyr0XyB2FUZM
d0wnoyYH8+mKtHBcJ7x5sjBuj17z84leixyLQrpNvNA1zmBL6zuva3y+5B1MoOME
/fLRiq/ZnaeMFjfWOj3ygq75Hv2eI0oNPdv+TE6l1ttA8LgtaWjvk3wE7rLUqs1r
2ad+h7/+NjkusJmDQeiD6ocfffEc6JWY6j5bc2BGya2ZE+BufN77NCtr3KZFnb0g
TEGMnuABz5ijMLz1PQYFKCUYlF92ZJd3PXCJrzaVoGrKLRdPs8Lq1kMyUmkFYY8h
T5TAFgWBk8Up10XVxNzqXjznzOPeRZKJQuilCsoT0RbBohQFJ7EVmL6Kzt8hR3oN
MwdW3K3OowstI4xhqse8zVrnnA99nfIkFiQ8f2B8qmaSVyjsDjrG/OrJxLYNbWBP
xMMY/WJfgZZlsIdO3bAA81480pgJJDNxrLtoQb71n8RC+hqkvTJ2UwJpB9bYjFQH
9mRmzevX4eHVEHDn+qs49pj8378Bhonpxgmh+XTld9RLr9RN64AppSoh/+vi15BN
v/vdGdrlt+9/vpvNRNetoyLxD/jyrAiGQEYCFr1QcPl056+3EgmoIo868Lof4R6n
bgw1mA3beuDysFL4dy1w6QR8fxxsV6OOZbOOUmU6oYgKejTEBL/Bdydg+wQt1/ZP
mQg9jmTDq4llxNXJcss+Jdyng/nWZ0yb0GI3GVj9Kgo3Vu/+KmmxAVxgu5ft4HKI
NQ+61oNLHTMuPEziEJ2m6WKFyAHOtQbeZXb16Ena8rTZ32RgaZSWSW4KDlv0p/03
pFTAH4tsDRMPlN7QesbDvVe3GQp2uhCNiUC47MiW6Ko0b45c5zGvBmYB/+19UFOg
7IsZQeAWghkMypsNaYmkWwA9DfwhPIQSDuSd4cFR4o4eD2okiUOZg1UjwdTjkwpI
YdnJKnMKsR1oOkota5M+iFgbHOde3bwAd/4QHYdUU4z90rMeMScppGFAGYPZw1d4
IEvIKobs8rAeSlr9YivS7RxgJQzZwu1E4t0B8E8kw2Sx7U6D+iUoBK7fnuDEFwhN
qhMsyXq6iJKrSGDQbwPyBmgWnOhQXafu7olXWpcRCYabrRf4xG16eh0HD7d//iie
FDuWD4rvH+NAc47/Oyjx6kwzLmtsSzgEzRtqgZZ/s+sbVt73UaRDUUptx19CuI/v
YVUWgXtaOm8GEBxTyGVNSZ7cHZAdFL+zvFiFfGYK8On69AksYIFO3BK+cFUWTfyw
jYmS/fme99OQYzXQrtcpwNElXQPPSH53ecETrje1tDEut7k6vZhLb4TS/K155abM
ditdr1+zAfcOGfl4XSQOD5ZAEDaoTOprVa57Ye7ZB+LQgbNwybcOZ3kSpe8CegDO
a9JyKgnRQ4WaHaUioqPjdHAtvKg5UUhq65sR95/cV6Byu2lcHIODZcUYMmMVLRX6
y7i6IzkIL8f/z94PmcJNMeQ52XwJDeGD7jaIhW1R5fhGLCPd5BBt8ct9fkvKpWAu
d7kGHbXKNH2dhyan6m560vOln3yLC/R9Uyn7G8jfVk1rbBZtzvpmgYXmCrwwlX8+
JgTHOuf4HDFGxG8LVAJgJphfujLRcIon46FLyCoTpqaTMvwRRdJGed26KD70l9gl
zEO7gzWIKTGh1eGcCO0Oku9Gng7nqf9u63F2AtD/sTOn1qRHrUI2I8U0DHitVpce
va0+prb/QQl3hA5eidj32Nfah/8tf2n2atnpuhOn/oGL3QkhLpPORVKs5OgqJLzi
q7GA6Q9SAyZ4yodHKHSzsRaedO1GHlxl/fAbkgcurNj/00aMuMxEpgaMaGbFhJmS
WtjDXqucO2QmiMyBhzXkgQsh25SNDjHxStTrsUF32HbY095U0TRZl9DTNNuyg11U
EA+M+YKidKcq+Imde4X5KbN4mSK7W6LYNJzio4oUVSx4AtKjhJgqI0ZEpc5OD1Dm
OkISC+Z/T6DS+tb2ABE1pcQC0b/N7fADShkKZ4UPEJS7/2SE5nZLKdbcEngh4qW0
Xv+AKfCiaOCOK8tiATIMOC2xhOxkCcf86tdZVTeM8lFwe0AuaNbmbKoQUkr/Q/2R
yossobV9zTpG1Kp0x6KbEn7SnHfmHfblPmS2HSmE0pE4yfpLd5lY7FQEsCMwJ4Wy
fPlbw+RUpkYxSzAvG5YBG3YHG0k2IynOzEakZ44wKOXUKgFJ/LTT4s1TbsfZhlV4
sbiDpcVhxL3JGVpwameHMbYCd4CBOMXWu3Kgv0mEf2ZOveDkjgfp1xqTXSfDspfG
NqIPGGx8qLcbsc4IU7bJdECawzvaO6NhlNKefUh7jJUEEBklxT1uIxYDHWicoO3A
4G7SobLRQoIdZoLxpuIWEYP/b71K2k5IWrIeAKk8bIOskRFnWSP6xd2OybresiYp
csHc/Cx4x+X+U59Vv1zQ3rjow671IYXlfUpcvehgVkK0iWH8wIjucWv6WCiJNYER
rI+gegisOAWH1pUWwtwQrb5wlNIKKbeABuejRtXbw6b1hoavU0yN2n/qKz5xDA8t
MMrSBFaHRVCIUI1/BsJO4mp+q7tCFPKTeqd60TciE8qAwW7FOIJ00uBVe+KIfLFm
/9bHDeMCMaOK31J2OwrSqFKWi94p3AT5sGYAxHSDxfh8IV7sONJKPUinIiLoXJ0x
IPZcfJo4JrZ/1tUdo2rZ/eJf4PfM2qu1dgMGzfDCD0C7Ghjp/93beWKh1942hmME
xvyE992+8ZrOXx/ftt5y4De8uc2Z2MDYd2x8DNjWrn0iYlfF5QLuzKOdkm57lszO
pT+V9c5G7bJk+NZVh5FJch1HZvXxQgvi8qXnkfeK499s5Ss7y0YJSkuE6IOH34ht
h7rX13l+4xJI/MgRLkWnLn6j21m0VPjEk5GnIi3vb+r7sS/fSOPHf87UPkpC1Lvn
+LUdHd1jhOBR/C6EEFGVlHLQy89Z1KwG0vT9n+736C6e3U7UHzDzBNL7eNudKvrH
+D6t6ooGocopdicqs5bDQe2Q9StOhVnCGuhBmSMkcpoQWV2oDy8wcLO++GQge3CE
qH6Sb5AnhMRZTPZzlDbQZHraEDLQbyFvMvo2t97V9T8MunENh/dmGo6rl2kHeV9E
PzPN2kvSNSfN30cr/tfVXwcjsrDAGWD52e46m5ZjhBHChup8I59/8Z53o8P66zo1
1JJLKIN9VPH//4otrrwpFlOCOssJB7Nc3oEcbU42htIXzVULZKwOFXlpppdS1pS7
YiQWcLY2WsJz1SdwR6Zf4bFOZfJK3ioOiIKjLZfrl3jdwXn0asxRZVxs7/oLPWOW
SGsLk8Y2rRCvBw+3v3s3kXdw2VixWqz1iEvIivydBTOTDBu5LA9OCxZPvSkGRDd0
EWe5Qlgjqs4wpiDhHkvh2A5S4ucCXtskJX6i9Fq1QVSB08asMo/Hr2VjRYtqfSNl
0Bn7VFSmbVomdelek0GPyqZzrdmc10zV7Xlb7YwcEbzu1wdyX6TUGmXB7opx6AfE
okSJNxLljdQJgcia2vtCjty0fJUB8u20bA2twV+nZpwm1DeZDyMsCB23ptGRb3ch
qfHcMJ8dLQ6xzghN+KWhkVEk4BNaPH0xXjwnkswvtjMY6ihcEsb2hpT4wFltXF8G
ltTT/XtlXwQj2d5fSe0VkXIoF/yreCAE27cLHGddE6Xe/u4F3YeVLCz3H+FcPyhI
PHVFzrwO8jCdeA3I4pQc7bG/hYenedhKpOkxF8ZvDoDar0z3SL5gdorHJQUtAA4U
ihNLoe9TrY3JgW3dXzQuuaEN7/eO8kn/We54lHeXt2ZbFg3KwW2KTkIv97CJtjfe
iowB1vQGT+4642Yev5Fk+d0HhFCwAXUmKHlks6AlqLG+/dBu+wp4PvLEOFt2GH3o
zMj1z4QPA1E+JNLbixhFXNgUbo0x69YfZGh/UCGgGzuoChdRzKHlGrDuldOJ0O2y
2Cv53mTaFh4Nt7E1MAAO9Jts8NEBLmtEvt3Z8Fu9iISiXHe1f+RA9SHUCr04wbE9
gcVkN7FPlKEf1siyLC22YAVjZ96af6T9bOeAWIgznXw5ThJusT9KbZWA9D88sV5M
WjTypbSurWayq8h1MgiYI9ePAZrQP1cYBstGE2FCJ9M7qDyXVri6jz5G7BENA9VZ
hXP+cr5qQ5wD9VpClv0SEvRboW/AWDPjYzemHQwLirHIPl8XRfsP1PHPLIgKkTbB
dj1pDE2KhB+APhyfuR+XDM0bYyo9O8BsRUtH9arSwJTSbzQoeS51MnmkuxOJgNtr
xY4n9HRITHBfvxZ0Qg/fR6OV9i0wI4WtRJSxq9GvRWWfkjEL3+02SdB2dcmdla9J
LY6TlL/cQ8GVYoy1BV5HXIVO8yUEu3ay6F3HyGex3a92nYr83lqBhsSjMNVw31uv
/gBC+dgkhlS1Lr65nrjeJRYUY+S+glGjyNXWhRdalrxCOGawi/29Lm5RGH/7oA9L
fg/Ggs5zP9oOZjeoKQavYyZZiQC0Obi7ydEPlXbguHWVAD1+SaoQe73zdi7Da0MQ
5P23nmEp6eXG2R0JlWY62NwAvr+ArdhQUQDsyZ9qo6Cu6xYLZjC9f6ZWUattrQ+g
erZa8cWg34ZZXzpARbIh6yJvkzlmxdp+JJYwJjT3pyqWzzT9l368NBHwqOOCqMbA
cN3idhpHYsqy53MVJGeK+8XTg0at/3+IZaAaOZjDC04RiUVWZFRpEEoPjbpDB1eT
/Jr72m1oPxLq/TxXOWTr5cnCD7R6sdvefevjMssH9EoHK1AthWqc2eNPjc2OY1M3
oy7zGuN7j9z3OI2HkteOQrODC9ay5/7uOpbPuGf23WZJ9r5IujJIrgRNMzSI9lsE
a9sy4cjHkeFFVQ9aNbpBJqX+uuG+/2p1htipck8B8plhmi9wG1PpzfUYqDP1I0jf
+XfyZe0xUMlUXGoBl11QWgi+h9ydof1XJgMMs/kYhAtqF3IcLzuAwC5MIpx+allb
av96VCUpDndhiQqy9TNL8HqKe3qz8eJgxvBW4jbwvwhtNUTOfpkWVstYLVeP12Lg
+HQrxP0DQ1B8JA73xH7NHwpj1dlMcrihsXLVMOUR0n+sAXiEUwLbQ31HZ9TVqzSr
qj1yr9ik1XXrFG0Et9dkOHRt+EhZenCN1QogsN+GLIXDPX/DEeIT17e8EvSRQxF7
TPc9Y4jUmtkF21DVnJstk8CwUW6bRAaCGG49FGMdpxXzLQw5+pm+/9y6QZ1593C5
qsaJUnaNJH/spm8OhzNZjtLH0wdIm0nrk8O0PwuNUpJbGUSLIeWEy1MKGCxOhlD5
LYKuD7qm/RNuh1u7swlX+AXeYzQNQ9cVZdhnEzfYc4Shi1rI6gLByrQmxH19UE4E
J1caunpLktRgJvRT0UirKl0rDxS4RigN2EdD0pF83Z30fMe6IjnDKnlr8Cv6g60G
Sw2iNRAPG8FAjrTjv+6kllMK+jE1kax8uB/uwaOjA94nacpfTLACH5UJXJg0C5NL
C7mnRDGmlIuXFcg71sxbj2ZIZwPvqbFk3gkxAINZVw8QHsZphcatdUuNS43h8BYs
3a2+09MWC54x5XHI/SRTRgA43kxwxb8yu8012tCfnVbqC8z5xnFxyuX3CV+f25pq
9aWAmKvvHEK8Pa31dNDn9Ig34+akfTcN9ZCzq3F8QzXWe5FngLben/NA8Y4nX7fk
rf0iUWrRTOWQhPNANfHHnTmvvT2g52FMAx9d5AcyIiMW9iQXGyNLTo23uEXzsQ36
7iY+swxJw5U2sWBf/W0QqymnHVsSyUQzL9GpEUqQOXSCCq6xF2RNEf43cAu2I8PL
yayQ5HTCet1cW17rxZCY2MvhSSFbM9J8tCW4WSjR0pveWY5QVQ3dzmwOEZQ9GWtt
oy5MAQdc5w8A0iCP3zoCrFuHS5iliHItf19pTxvGtJBUig+F/YW01Y6gbfEtkwLL
9CFWmxiPeU4KSL5hVjQEApguRQcu1l1y/n0BvTNAfFKHTmsUEcswlvZeG2Des2wK
MwZJiTudtiJ5LJE2rNH+8XrqryRI1+vhyzuAae0anutRKsCgTVSo3SURWdqisxDX
SWwIwRLRyUU5+M1oHXP4wDMzHwsgfMgkoV/4eRed8MpGN6DZC1GCXyb8Cpg3Wmax
LMu28dYQMuMnZL66MgQXtQj2nDRjbIk0sMGqvD1CDMuXQUWV6+/RhqPxZ3tBU9jD
YC1PMmlaknw/8o8lY3y/7zas1OPDuQWD9+quABWucsK/atUuZGvOdybNtg4Y9rCL
nm+U7H2+7yTXiV+4EMjRtxC5ysGC4IQGYuEq8VwYvMaHSlQ2LvsbJ7KInz8dlR1K
sSXn7GBfw8dnkIS+iHikwjLRk3DVrbY2oQpQWzg9xfuNf6LWD9InglliPQ3xoXkH
64ibCWr1bTtcqnD+bqoLbZ+E9LR29JlXFwZwJ2dvXBAOq5erZiptJej968VWnLkg
lmYxkng6EMJaqjiSkewdzMRSzbuRGeCbFEY7WQeK4nm+2Ckn91TWLuOajV6WdDzX
+T57Ctx4VwDO4cfCNv1+j1idB8wW34AmhEaG6e17s03xRNiQo2Rc3ipzlhAQcpAC
1A65RcrIv7LAo78iQk2Y8VYxJQa1Qn/ugYaNtHAUFg89lXRf5cxBRd/tkWkcBBh3
XLtxjovHctnWyk/sLTdoIK/PiuGUYs/yw5r60ec1MV3hHVBaX3vVhkLRzUHANTut
HUAUibe6y7hAGbLFQjpluTAXDPpbKQsrLL2/BH5LKIdmyHKFtfAk6GM5fd4I4B+N
BJdfucFucZqlYCrtWFAvaBCIHs2X9PBK+C/IKvxE7EnXxCe+Lj9pKpHKyMmB6oaV
OVZvRPfrYCAjQ4Lo9daEHipZtTaeswCtJfgJLxBQ/Szjcu96z4akaNjNKjn/chDE
MkDSWMykU+pHM4+Ed1oGgByjEQ84gRs49tOtrYBbixviUKw1MQWctuMv0iQHHOfF
HgsSfghJrbDk4A5SC6zBd0KzG+7uo0ifCPErKZbWSeAbx4r0J9HtM7XVbbGTSqnL
MCJysYj5QexxAIUsEWaAc7GHomHyD3SwkbYpTBDgphHt/iWrESZAQB/qS1FkFLc7
OBnrdMxwaARUEwje0HdlDCprnjOIeVslRkM+v/xOgvyasV256aOefy8X+a9uE8xP
ZWb4wWhUTpaDyAJ3PkIiBjUY0I7Fy9fmjexjeWzcOX+2Afw6m6cg/feJFkVaHKmv
hWv9p+1AssKilkmCcotGMbQdXQQqdeZK5qgL3l63i4tc9kAmQL4aavCBjC+jceCJ
1YnJM8C8Q/kV0NxkhjZvxA7/TSt8Inbw9lLeD92s8nZIhbGQip8KDOxVdRgR3L8C
j2+ws/MrQe5U3x3SV9NbsJqr8U68Pgs1wdvGO4fpozcn3jlZl60SGvCa2VW1gcpv
2OCSh84SdTTXQmViattRquXyc0g4BQ7VXlBHVqafGXqMVq8LqyJM/jWOuCVqRXSk
mzPd9VdEjrOXUGa3SW6j/g5Dy3faJ5Y6fwqII8hYkXT9P7fff22f6WDp/IVicOAw
l+f2T9yXTNaXLmVj1cq6RRdq1UteQqE7Ts3yl7Zckp1ljJygGlnbamYifu5ypZ/y
Dn/d0V0fGQwpyqZGFxsSzYuwUqRV05TzWeCeH2YQjn9kRtx6hhT6GgwBfP1bcQdx
aJFwAjd+bD3M2mMLzBp4fau9F0Vs/JE7TQpL0MRt5ofY1iNiLErMkTx5KwBA8G0c
H3oQ6hX4KaL6ERyR72F1dPHNpfvL1F1oFhtzvoBv4RdB33kpjfvPEPy+yIR25JgG
EPV6AceR7wiUv2P582PrXJF1VkruayIUV2BR9Tico6EqXYlv46GKBFeT3q6wLnQ8
SMbGY894PfIIE4padybGbcP3KMgC5Eg3o0sN7Tb+dFRu65LBfCoGnLMKfIpAcvOs
b9QNQfgSmaVtkjbaxI+IulNb/eDeN2HWYU4OeaOPqGzlZ5gL2T5nKSnFYLqTQ0F2
9Ys+LMHGWfPgLjYP0tVjOEkYSjhxulW/T4+N7V2YiFKMD2EeYIgKzpwlT4k2BsuZ
r8YtuG62j4ufjfiEeOpi4NUPi0HpeLRYxp0HCoHvvBvPxZ3rC0KoU21FBDOVBdJ6
1m/orWUK9qof2eBVbpzqCAf0V12lgLRQ2sRQJy4+RolKDERjw6a+EImR1Soqhu/P
IJmxlmANOGM81J2YBA/ieLmrtU5uLNDuQzIyjbYT7CRGkoDn/pDhU4JVQWRbjkvr
OlkW4HvE1lpZGkVHN/fkLOkS+CNAuh9X0vqXcaiBCUHS+kfUoVyzsXwpdnNflp0r
XgvjvDWLeN3ld0L9nGT1NCwYPfJ1ExDE0HHtDiCcOlICAdTmXSj0SpQfKZvFV+EE
zWDoNGD3WSLhQG4gOvLr3xGCHJ9N94m7Tda5WjiEpfJOCiAsAadkRryo5TFNm4pq
xOf7pLj6armS5hF5DgrfQRx/5QbhZqSJLHHBz8380dyqpWYMeGlFkQSqfw74awaj
ZMplyCjPaqGZ9DX3mei8XYHyqNnulroT7oOViBNkcUniPjbwHWOvi0bSJVk7yjYH
C1yL07ss0ztuQqATs5CGSuwjqF0DnCAnavKNt0WziX8mQXHD89S3MidViNKMXf00
Jz4iiBHsiYuZ+m5u6QAGyOWrkhGDQaWQlx533y/yHgcSgxZxs71wqBJb2xVFVLhg
SY1YEkbT2XHNcVOxXJ0KdEArEob80jIk6aujbQK1Z4p02ag9a5/JVknFV6csSIgK
fP7Bjw8YU8foaMKI/0KCaCoWmeEiIb8YyWcOfZ7z/L46q3m5buyYLjUbTiJHCu9j
wryYZdE8BXPTPta7NfPF9gp9QKv47SBf6BYU25/3qr/bIJmyOmEklOR4M9KnBZpD
jwEjqBuzELJ7GamZx7Shh8NJQLD6NYzYaH1o80hPN/sJRuMXvwxACg4a8wNB5dYS
+y18JKKEhmVLR2A9tp1xqlidczgVcyaVJ7Y40HAF/rybXZcUZGGn9/Hm0SvvrBMq
oyTZ39cqx+/ZzA0TwVsGLyqPEmyW+Eoo426DsUYXz1IWEobHfr4yDxG4Bb/hj7L6
YXo/nWPV9T3wumSBW585QIIhCar1Gk60iAQoUJlMNohUuj3F/hiZtVqwKsI3+h0n
R8f5bdr3GJfw3syO4w5jeJC5Q93yItPQrOUrQJuBNCZlaInG/Uc3ZaQceKEa67eA
RkB8wPp1U3ba1gxoz3d8JEEJNdZtvjVoRuZtz5tj2oTsw/jbUzkjLudyxEX7oRdz
l9KE5peXQAR0DKAnoOJinZWbFbesyHjiuNLjOGk6+D2VIndI+x7Ie950I1cWiKB+
J0MR0dBS6Cczl7hT5rUR1yNow1Svpd3ItKeGYPVuNLFKiATccHgFZjW3CJ6pRsD6
5knHfboR79IKzTQHvEg8BkXRBFaA6BjX2dEK0k61u6xbvwPJTEizPh963s6OKnom
PXALMO6oXY6L1ApbK8xDaw8Xfu6p7U/uZ2WtphjvWYxK1qrnANn9R+qH3J6jP981
EdMIdM+rsy0beWnGBD7b+bSFA+arsVczBoUp9E1Qq0oHn7hUKBX7ayL568soC2aR
Ot6REyEAISc6b650fisUjLGhWiayTwdp4xexiSkPJ9Bw7ngVeyEi5Fs74y5i+/Sp
Bl7uQYBw6CIVYbKJnlF9lGK5+E5CuwA6vZUtBcyxXaM0UEDNKVFfI9EBdZduCrOD
pkbMGoP+M1iU/TApwo+qQSVDngtyGJBd1wYcceRZn8D4q+A09ArpFNVdXDHEEoj3
EE7/Y25wLqH+diTVj6iukzWOaXF9VWmxnG1yxpGrKobhn/gfINdyL0vz/dbD8ZVw
BgybumxW+ZVZaREQ3j5r14/uNJ1pAPQZ1rzkjNnBeS/7sIlAdz1eiVg6bZKXBH08
Qs8kIx/HAZvlrnZRbiN/e7OQ11STogM/1LTsh5JQa+38xMBlbgmc6J4PyVZc4pzM
NeVCwR7Xjb3XCsmuh/CoKmaZoGiqWfyX4lidzDnE3H8pcfjayAet3ZWQsqbfzFLZ
rZnykj2gBg0tbo6SNtqd8SUNL8OYm90bdXcTcpOBZZunX2UbqtEkh0Fy64JTNXck
wfpuB2FSk1SfjhD93V6txRepvuBIrPiedUfDJEIgg9ANnu8v6Hs3oZjrfSC4S/MJ
GBgUQqMo1bo44/wq54iBVh9CpihW2CngB1HfdOUDKSxCGRh4eb6/mW9UBLVN8SBt
y0nV5inJnw7Mo931cyWlmnR7qfjb7tEbkV9wFvfUufADpNnPBrf//UBU2G2D7RP2
bf9gsMaWa/q0B70HLwsEatzchTIpWXN2Icp0FjW6vmoNR2GEAUTVkhb/WM5Z3EFp
xldt1RxQhSOKVt3oHpZ55y47vJSs980A2IwKIthir1H49j80hXb6VctyZczwxCWB
aa8I48rv9DdhI3r1nwT4mFKMhU+6cS4lnMT784uS7nF54CuFdqFjsw1NPKo1+BcF
VFe4cGv9xiwUe++6uuFHd082lOGfu0gywTLvj0OxPnR4tv68yhX8SWUx20DuR/lh
IOFxDBZGGoaX4jVvs97nlmc6HRMz5eWOwX2i/4+KLqguj4RLM87iaFxWcilCp/j2
+UqDXWc/v4XoPhQgVraXZUH6wWOLl4J2M5oaZBtMPplJWvbgb2yYD9f7/0yeKrm5
5fToC9KZxDH7jv9eogYpMLLeT3+V/TrDS/ax+F0s7uLe3JEf6bVzIWuyAXMybUSr
JDFjHLmuZxhZTS6qzfrPe26i9rSJLJVMUeIXQ2etqTl9SwO2VYEYFLb/7SWNoo4C
QjVbhQfCLpGOQXn+OoGTJVRU6KAql0PT/nqYw3rRIGBx744LaqMZIPm4ltfg7Jse
7n40j/ojrfWswQvjaBHh2/rWG6sSCWEj6q5HknguPt6RFJhfjIxu9LBK/M3DkhBK
BBPrWpYGn5b9r+mTfR7DFe6Vl6ua4oDECL0X/hyCUw/UBqhsXXkH47Q07KLwzB87
dNcXI5PnxFjZQX4A504ERcovg6VPQ9m35tkT3flrNmzQcvh+hvbpqaPT4K6uR6S+
NyuMl21cUWuxu80mysea/tgLgGFtfnrGN8edqOam5Ma6XDQgGy4IUvVnDWR+kve8
UgjwBnQGi8bfsykxDhmFmAJcM8IiTsxmwSTy3l1OoxmkhHRvG3TjMFnKwZtdrA27
DqfedAgWywe+G96MYoVbbwWKJnomX0vGbBUQhS4ngdX/DEm31rA5KNr9ZEtGjNDe
rOsrkJ65OgZXaYg/5nbGU4mbQ4Ut5p7/lEkYGawXzPQOpBvvL2KRkEzBw2oBtoKn
1cbx8o1GfQ7a9SBEVh1P+jC7V+TBhmS5Ux63xtBTIMPYV9oo9i14z7Wb+GyUwbuS
b8GyijthAMKtB+h/iipDxFkO4bigAE3AHeCWdM45fwI5F7uJp1lRRUmP4fHJZxP1
qCdPj5+uhhEQtDbR+XmOPuFlXu0UqXn9Dl4RTTXgtMSsnfeiO+FJ+npvk3t3IWSr
8KZ1OiBusowndudoQCg+xYd7Hh6MFpEOXnnXGgtMZ50604YQwhuYjnFM4jE+9A/u
nGiD0yek3yNlZwPdlfoKiehTCjNhnGrmQMNtq+MGTF91LYORkj4qzPPP06ZcOXKu
f6WE0PVLFCIq1GV7DoA8i05C9QNRdWvGSZ98PvmifARat1nLc7yysNriiB0EMXzP
2qOjLDh7Ys9V555lfbbMgm82BWEWKEtkELbD0jq4HR/4DlQ74T96TkdH3upyEwMs
ZELuec/vXTGZFVLsMwaPdNzf1DTKO8gP6uAcmOj8ffo9X+FLLcFDKuyL2xajs4fT
cs02B9/Q7OLw6g+nrmMsNvXDrENQVhLi2FlxWSKdw0xmJQWmMXsYjHhi18l/rrTh
3veqpBgjYnzmOIl1PyUw4dsCYEhTDW+zIjMDkMHpk7VGXQ85onG84kGdpveRpNE0
NiYhMztJqWmKZH5Zp0Rk+49b5RAniFl4IyLxXSykQHQ9DAFL/JW7QmYhZI1+p3Tj
kypyKEXewGimXaRL1OSK8j/0md/rIDmMbkzHHxfbdu10wtNNjkldunyLOm86Rnez
UFcYlHeN6MfsEFcYS6M5biVZniLi+xzqfd9AoMmgMSLB/ekqSOn+2D4M+ncuqL8+
vHqpozEpgS9mqRMVksYHhsj4b0bMWYLRUJqoQxPn6ZubMPQ4lDpUNt4FAvLZFV5x
krrITU62cg+9IVMHd0qWzMqsk24uxHBDKSqD+f7RHUjdHwlsbnsICdgEPKjf8ucw
TL2kzVlctoNzIi/AjhukPp6NcaAj46TFCLYpJ/7pQiUhYXwIdaZPFoYS8uNwG2xI
nm0GlZo6xNT8F3b9BP2/7NbB4HYsvcC3C0pmvUjYGhwQKdk9qHDONtQUsaS/IaBK
gRSEoU0pQ/GSTZffL0fx9aYztZ021hOH+8lwWPF17F6iRP5QECzjGD2+Id6LBM5h
6um7gyQiY3fSY6oLUA+fZzEh8gfo9NzHsWtAvfHRj7rA+4Wtgq6RrDshp4zVbfH7
9p9j1qoBO7VsZFbgPKZD6Uosj4D8UDIc0mWgeiTUmUvEF8Q46flzMfz5k0YBXYde
MvC/92yvY9cTmU3eflsZNDYB8ZGrmznVl7NF4l69b98BXw8rGqSoxrT8uXcL22UA
3XB9C4uoyd9CSbU9+QKO+MDcr6NLPg75WSL/2sJ2wsndovKxbVbNby4bUuTEYtI3
vDhyLp0yHDccjxvGoZCxWwzqiQCZDXKANvbl2cNQn9HgzQAds5FB2XHWqkWyRcc2
/7xloSKTcfaUCoJ8my4s8/vn7Jp9t5G8Vx15W/dkwsOWQfXIchH3yl+W/V6F+u7H
ahk7ipoOptFz4xLOWJozx0m7lZlq/lOpxvWhmfOc7tbrXiqLGxjLXU97aTwq5sH1
qtlhNGk7gdOpNIrQcTGPWFjXwCUnYKEqMGf61UDSCt2vt8UKQFLT2Gs63ENe86t3
u0Oe4LrTRaZk/vXfe9Y+kQw0HQPdM1mrG3yrx4hBzekZO78Tii/SNsaKhBvFQg/B
60cSRCYlYAjsdOIuhw9DTi9Gk52AY2O52LATmPzpXJ1vQ3/Wt9KqMiswIs6hruzc
ZnNsyriuRzdqvBkNx99epy1fIXaVp4uz/L7xs9QnA8VhTY42V1Y1DYbjQkwDe6wm
wckB4KF8weD/IBlPL8xNc4oD8njJB3fZ5ui8sJWWgfXvaAkseaxZ+wCA6UC9Th7w
jCJ1mFMs22/VpAOMpn6FNd3ubcjRdr0uzvz0luiAIuIUGbqqxUOfeV712XfTOKNl
NkHIzXQautxcuDqze7vD+daD00icmHhFSm9Tm4BD8jauNrYUWhoHKUgAC/I0Oe5f
ykl+OJcyyZVULN1UDZUOOEfa2F7+pJ+0xQkx6dZI4gKMuB8ZPRAp7ANE0ztW5ka+
wGOS4+V9hRrYEtsMBg7nC7TPmwQtzX/v/FInrIRgaUvlfNOql6T6zbbzvXz+0N2H
6z8nvz6fJFVLiJ1n/QaoPraRanUxk05uq2wZCPYZ/n/+qq5sSZUzojChENwcNi0l
+6v+ojsvfmAsq0SNc+vkQeECEwH6TMGstqDUkmzD3KzO9XkXWS3DJ4XTYYbhcNIJ
/YX3traLEyx9joAHj5x2jBrs63NAVlV9SZTBu/l+YYZN0Uz3soZwiWdewTD+uFxw
lV32fd5PaSONiSVoXQYzy7KW7mJG36FYTTO1I+zzMXxoSGZRCbRpm7h9xLpG+hEx
einHQjdQ43virIPoy6zYk1QX5hgeMJ7Z9vNRZY0R236YWdyudPqc3B4a8XJU7rgs
ZJuqwMR+szxvNlFJnNIq0iqo2tDZOtr41FexuAehokbLA9Y+LMQ4Xmqj/Iby0nUN
KruEzU6Cr/u9p6nYyXtRLhFVtkw9ZBRa+yJLcgjfLAVeTq9yTCPDlJAHoNWWLXZl
`pragma protect end_protected
