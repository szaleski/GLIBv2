alt_cv_issp_inst : alt_cv_issp PORT MAP (
		probe	 => probe_sig,
		source_clk	 => source_clk_sig,
		source_ena	 => source_ena_sig,
		source	 => source_sig
	);
