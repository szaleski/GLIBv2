// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:47 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
XyMrNCkkvhNKx3gSkAo6VPjYugkecPM18i31JC4Qofg1NobvTezAOLAmAqJ2nvdR
QGu6Tkx95/mdPtJAV39y4MAiYlX1G8NbM9HwcF4qNBQjBbnQThFBZ3/mBLYj8aYY
gf3XcPa0act6boceHdULNAiePtlK4a75I5j2+jzlhFY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3632)
fl0n/GPjUYrZww2majmDcQuAWpsvPtU53pqn16dVMr+JRnLrkn+F8WyY3apW8o2x
skohRotoXEKwHKoLY3ZHlD81C9FSZHR2EHFLKAIf7tAgjupZvHRGK6zku2T3LWcW
GfPfBE1Lwl1FZZ3K20iIkBzv/C2Jj2jiHYHzMtEPrzhM2IGGcpO5fnjSrVg748y1
MuN2ZB1xUEPK5y5vxbiPX8KSLeeRmn/lb9Gbwr6Mgu1ulem3yDPtW96U9nVKtp0n
43xu3wXxiM1QBxFnlIGAR4c0ofU3cWK2DJmFxHgryfx5zj2Uz14WUBKALtxlz1eo
pX1iHkyPcRPr2x+lAk2oMNy0V0jlklu50RvhGg+lqsnmTD9SN+6d/yJMAfrGHgeX
wRhOHCuBeMYPigI5BHB45n2+w3sZ4UOyqQC6FPpBeY9gJ3KQuEzgMEC5XnW33xCg
VhAsvVOP6b82KFaQFWDciNk0baXnig0cNZSdEQLjmVhkUjx09YffijIfdZQg+ryC
0wXWCnTkI0g2TXNF9HYmwSzkkraPWpkv6e0K/uEqyaMa58ZtxS/D0HU4kaStYj5I
2V79+nRV7hjcLEjPVfFGZ9I8NoAILWM2A0Ha3iP/ph4xNmdyf+gZ6OJlgABoP9yQ
DSdrwXUAS79CapuPtYW39Qsj0R3e81jaObTRV59GFRvTwWz7rdPJcVOdN/ZZmVLZ
N5zHrhs4NwtFOjv1J4yWI8etblSIflMztrRry/BsWJ0vyYEdPiYwPdgAgNNL7YRI
HzbWjhEjIHejrHllUl8S/IQQ3NtqGuQ2Lm3S6nqx08AwerFMEsc9sQo81Iv30rss
Uk6auulsImA6QedmoT2VeuHoflZZcQzk+SDeae2XIB1f9esfkgxBI8wzcFyOaW67
kvYMO1iWHPK+m8ThAs5n3R4YNwdpj9TU/FqUHyQW4DSBFrcixqKnQbjzfXL6iArK
z8NFGaIlF4GsjM1kDAfaZ8xOot6ESSft3YrsAHTYmzRkPAuhYJZ1iwf6zAkYVXDe
2JyWFTfj0hP3Ob8UxI2pIMNAi7r39Vf2NPKst/O+SOfItOgM/pRgTsHXs+HiIfRS
a9YoHAwGen3RfXYtlqTdER/2JLetMMfSmdR7CIAPM6Lm+iKgM1jQiTPnBnkET7hN
x5C0VliXQPiF1s3C1bYHQ0Uvfpb8BhyyVArXvsCE+Mj91rnqxi2Mz7NKCgFwpRZW
mTXtTf+JSYOkAo/7c/hCCk8vvCdE83EVJIHsl2j+P+1WBxJIQCZFCU7cuT/ntUVg
NXj/pxIZKHfcLgYumZB07ONlXxqX5NEjrrv7ndC6SVOA0ANY1/mTJLSiZu6r6e86
NkK3cYaObxvsJYH5ZTmeMaVRrEByl6yhNWwXjZYuzPd5V4hwnFlJO8YKiBfYo8ph
259plW83WJxB8glAR+wdbH+GS1Swh84P3EsetvyXI32p/RhfphxZhTk81Ga+tjbL
nFpltcI/k4JNZd5xEkBTJiOvI+rfkSJruI7DPq5ZqA0W2LRGx/PbW/fY9aQ4GQHN
Yp51OWaioP75SyJA1MT+lXvFPNrHyRviHiAIJT5XKzHbPrg/q0mFeC3DvwDt4m3q
ltWG7P1tPG5e4ZTGej3i8IbMVXda/NjZYhP0Fb2mi7zEWtVWo4mjzQjdk8Gusd71
2k5ECeqpDUG/vFKijCE2xTV62YRn5Z0t3cbI+NHO2nMHZMjBgLrpy+YGREFDI2d5
bnuLHJNuRw201S/tGIp1EGAIL8FZSCvTX0qsoVFkUCVIv7VnFHgLeWTB/3QADhZ1
oQTSVuyGgdZVlFYBE9LPpC/0odltHS4WfG1bcUTIJ0a2C/tPyudzkbZ8G4K0xYYp
FttNY4fPajMfpNI71SaJm4nY8Rs57pgU87+6Yig/JXjcMeHtrFWaW5ZOxU/0jiKz
T4idLJ0/8DNrz94uKn5y16B7Or+r1g7CnrZZmReySHhf399rNnJaFKxOwQhzsPL3
q3TRG5BE2r3RjKJjnXe4bo87pVlzfiVrNCNy0wmPW69oaTQpzZpxaECKPGPDGhmp
Y3OEBxsyhXtejb55DnUhQAGbZ+1p08GjB6p4fTLzlcASk2Wn+XPd5ThjrSfZjNaq
jREiotPCTRxtLsGET0iHekNj7BNdwOGWtjmnjjBog3S3R0Vx5LhYbZsUuqeUCwON
QaAiMpbh8HeTOnlC3ydoBFBlBWc3P1kbVK24gRO83f4YDelrrti6LN2zXGB9avLW
e20nRv6mfgkqVugM4WBHQOOAhuGn4hEPHkVhl+9syprahw1VhDDgZXzXgXk6dgLc
2c/aisfRP+Th13lZcTeK+kjXIKx3M+D2k0wJ7oQuxPWMAREwtGvwEuucKuIWnXuv
t35eBM/mVw5oaGyqmQfDb/m5UNRCpZKX1cPiyfCuQJlfmQikGb2gGveCVROvmCxS
dq2+RjH92hHTliZsFmIjOIj5nDnLlj+D6YmgSD0gF8riy1hjE/SmvlumrNQBuiFb
EQI/h4sRJVzPcO8kjPgC9mAWzuC2zcyiyvsi2a08pp9o11o16sKlT8x7v+ZOKM/J
D3lZNb8t8QX7xGQhPhR9gKoYZ9T84QGfv0BjfQjEyBrP28f9iR6sQ2Ls1TfMswOC
jS2lLBtsQ0cP2jCIi3EF8L+WEPsQHZlxYGgwA9R/at4iRfoyizebSrC3gR+XepuY
bDQg5uvdixtaPbr8ekSVAb/GJmI9l3rFWpxMY/kZzvRirPnjU3gkp8+erIf0VXiD
tvh6S9K5PHmRXwg4HyT6CNX839QDN540a+trvaEpnNeqBwv3B/T/pqIeHi+CIfYZ
KDQmfobL0FCR48CBTPtu4K6VGM9Ia0C19cFI1KYqrplXH7cMjFG1OqwervcXUYIT
vwbmya4gcse6Pj8dRyOc1p+OQvQWPet9mT1t3fB7gblQ/PxaP7MhnETac8cf5Ptg
l1GQhv0+My6GjvJfugqlzk+AWY3oFXWcgdROeh0YDo+bkoXGFZENOXWx1Mf4Gg2l
S8hzJQNQPDqWfzmJAbJAfSumFPaZ1OF8HmTXA4iUuXhC+Qp7tNzWKBlmY3X8WWXf
r9OmiuJy3ItadC15g0OF2aNnlWqp29F2EPPE2upr8euHVEGi5o3CaeEK3ybfA1Xu
Fjg3z+UXUy46REwnq8MLE5cmQrjex3VocUQISCX9bXPqMJPZ/jE7UimASFxEsOus
eqjLw9RNMi4kLrfwpHCJJxvk9QHsZHnNARgdD0z/qT+W6ORQAXvCkjT17FAok4UE
E+u7AQuXeDUCPzBuzQSuQ98CU0jXR+6XH5Azd4oJ77iwDSmtCLRflbO0+c6HQMi2
3LLUGf+TnoDij7Dc+UJP+jL6dHtAOBQ9RwVeznEA2UX8yT5AQwBqCq+EWsU0sGMo
XzR5eJPbEctqYQxya/hF1fwL6QQ73Ff3yTtFjBPhwsF8F8kpFcH2TyGKW8DNbKyg
evyBXHglbYvy5BjlPwuAWs2SxvekGVQ56a/Gd3L5+QfB+8UVnjJg4FBPLhpWlEaM
Uafsz4/RJs/xjT9z97sczzQFw+7qEJrZwX6xkSR1vWrLFNUvoV6zfC3iFG0XN3gk
VYdeKpAn4yLUVVaIYj/EPmgm6X5w2PLI2lVil7PWW21T6NNmp/03aC3ymZ+ghAgx
F6SMZ1gFvkMUbEB4oQ8UrUVcRgRazd8TAwiLmJmA4D6VkcUvC6pg59wvt54G0XaB
vqV+m+W8/0pN360Y2vYUyeqtlV+aN1s4pcvDQOxZgGOwe4vN0jarWebdQpCQpzpC
8y+Bp/Y03A6oHlmoDZYaz5ZagVFlvqFPdut7Oyt6Mez89jAsIm9yfu5QWVTjDd8r
R+sVI9pAYBiSCDys2UU2qaX+2ocg7V1X7T4H4rEPEbiL4Lnubm0rWG0UOlRJZ8Ln
E6vwSHi3DSd29U8vuZynSAadpggnEHFmMhiO4IlwFAt0vK+U0Kr54TzSzupPlQ3x
/qHuV0FQkLKWtxMzIXZVSj7W0CYtzRl0Req1kGEr2V5h+JGwheTEr37GuiLOicMT
1ActHxaZHkuEaMk2eqbVbiio0wJAijCpb+fgmShLEDNmvqnUrkZCpASjlcI13eqM
86+4CJ92yATtX4wWtb12oq8OQd4BuKTLSTOffuO2jestNB+94aKGMShkQekZAJg8
GNQhyIlVf7+MC1fh7PYJYjWsCRskmmgiMy1rvrNDMl++CR+uY3RKW+yyd49sWaq3
PGlHvsx0qfuQLqJxVZbDabv926HlMN1ETu0BP3fgcSrbWk2/SIDtSKW06yQmoMp0
MNkbsT3srRU9mJqROPUhyiuhqL5VTjMMmKlbRb453Z0yJmUSYW0kpufRVzLCGhkM
ppo7sRMxzIgXnVMBP1/csuGncrsiV2MFB1Khqqr4z8x1+Il/PwkEwfu+BU6/UDlQ
KB/MR4Q6+5Cp81vAAMbSdxm+dUjboYYLTvERuClTw0G/CsXj+OCKvT/ZAeOjp7jw
Qe59wSzI1E6UzXEwewPFGTNI+oqQbom8yNP199Xit9D6xONGhAw/gatwhmkdX6Ao
+nze1Dx1YwASvXWyyqx4vHTFVtsC7YODeCbe2uQa9eR8hLv1IdUYCU6lg5UyZLcP
XLbmkkIiy98C0pcnudE/z/4QJz436BIcx5Gxieizs7aaYnk/VIv7TLh5Rh/tsWlr
IyWGaWkgocVvM/LIg1vseT2b4V5Y66N1xm3ZQl6hy3F9LQUIjnlHEXBhG3HZkJj2
cpQc0iDDImP68fkUgkYZ9I8BQupYPPEwzdcvvUK9cimXRtH3aT+CvUVfJct7u0ov
aclKowA1dwbqpnUWS4g6JlduYN/9h10tAVQKdfBsv4o=
`pragma protect end_protected
