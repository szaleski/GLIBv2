// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:48 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
DmNh0LluaRdN5VdVayRHkQpo7zZBaQbw51mn1fUO/ttJk9OSB+LowSImeR51WyrJ
DhNGUcFNbC53cqU+GimZ5Y/hnJqAJISecYgSsSNA1h/oVAT2eumLw9RiNgLNMoS2
Q0PT8M0atexjpmiPjKxmkbyc3qd7dR0dH4HlzT/vF00=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5408)
Wqs5eFj0n6cBI0ggCy1vaXy/Ayyqu6Fc+X1cOfSbUE7/99r7u8uam1akYrA0oDrk
RXbIEPFtE0T55JZG1CfWHDabQ/4ln7BhikMeTXcQPHjULC8/QePrXSYMZp7f6Ugd
abICdpuhsZMIH3o6mJ4B+h+W7pwS4nzUwYKmv68vTtV4PSloJvkAqQyNftYr+l+i
W45wupZWPDk93XmkE0q5qZ4kh1FIZ0Gl2jp8ZtKMe6a0cQUbwhxYAavmSPxn+e5N
7sf0llgYzf92xdLrdzX86XnMHBbyYkVMf2KM+ZK1TbYphplN8xvU+74uenuKWZkE
GnCsgJZWRDrQc0IbOj+ZOgF9RLVTNpSETfrURPDd2litnPRpfZA+xUPwlO5nvOKG
fhgQyb/gtFRGhMSxhY2zrE83V9AfNU2nwKZ4IyjhJaQ8PQSrh+1i+obl//pxvxQ+
sO3vRjR2mv5xhEqvbidCLWQxYTBKI1of1pDMZigggpBGE/UV0UJOQeNMkc3Aq2cf
SzJkbImoGhVsxvNjWLIJhqJXyD+m49ffNNHDYgUI0+TqC0GzNb1IjdGwHIfMVatd
qQKJbXExz2qJuspMI10SrgaaUyeTnG43UVUycZ8LOgvtAwcfMHf1/Q84VSTkpe20
WHs9yzuQSY4pJKS3yg39lhUnSyj6EASZkQq7atnC3kYQs4/VIJdrp7mNmNJn+bn7
vkIefGdMars0z7NSVTojuoxHMBejP2Cevieg6NAgxqv+crOZMRIe15AQrRqWzs0U
HlJtsbROE80b9aYOrsfp7NSQpgP8s+gUErVn8XnDqTCLp5JftZEQjwXQdEQ8lhxp
v2w80jLjfiE5V1BUG0SNN4x24shyHyWDN06UD6h23B9UjRihBr7LC3jetq75XQ+W
xPTRz0nN2X1ESTn2jJUuLwPGrTWoCBcdQbSL0I7oTVABC4amoY6Yd5uF4pQFEUX9
d30joM1lcTlr+CbDVVV2nsOscxPcHhGQxR4GPpIwiPieOQm/q4K/w5Do6ivgUAVp
r9LrVmGkHOiYbe68KPYZXibXEC9ez5ZTvJMU23uN0IOv9/pcJImodgAtSOQnDwA+
/OpME1oHua2XaTPPcOexPWfthR1rB9zM+xk73db8h0puT0N2dUohUK0YfjS5AVZy
Kse9DGMyhD/B97IaUxm1mwCJL9mmJ/1ysXV6hIGKFbAMExkxBNLnxOLkcazUVEC/
xJLUYv67aW7QHDRXGna1IF685tc8Pr5A+hczwuGTEdoCoO9m/HoDnd13HOpKmux3
VSzqM+K8rPZknLLA+pkqf3022JvW8DPgJZcRVdP1LmA0dCOcUu89aTjOwD/hwJ6i
Xru92N764VvaC/iBFWgtJ+yXWtHyBqh7cLFwZxPtqR0LNVDsDyvQy0O09ci4AxmH
59UftNXI6hJVWcVPFJSEV4kVKck3ZTqJT59QpCzaJ9OSPOxIFB62B/kSGEKsl19J
WbhZ7XYITR20L7fBGmM0mJEbxqaTE45lYzVRuvm6qc88M9TIYwdWdAzLGfkzJLQp
2Ms+an7OGj5J407S2Sjd4paMpQUffTBPxsvO3X1xiq248pU4ezDREuHVXia/IaG4
YyUCOaD31M/7fk1Qb85+Zm8U3yiz2AJ9508/HyZLJ3jjEz7txLUAOu8ijIHtVT5+
mUd/v84BM6GIzWPIWUiSXZhQWmDELjjoCr2aN1oBSRZPbFGN6PS/xPfYcUTiI7AI
zwofm56o+7x7P8ZJOOrpTd5cLU8AQ1aS6mb9ZE6q5lEz1isa80k5+yw6wiPh5Frq
8Nfp4YDPLyzUAzJGQmhgn3ufnuyObUB1gVcE7+Oz3arczT/0lSlshK24XtHbGotz
URwF+x32SafdaNgLfHYefW/YJ+aHxSI6gCN83BApg3bv6gN67QkDIguEsC7DnGqk
BtsFH5dih+XexR1csres3RBYDdfJEZ3LzvwFsiqutkzspLTzcYdd8JCVEzi1cfSS
lCgJP+/510RJ7e9RJXBNKReZe0LFIFQjEkwPpAFat6ZvofCTih2kLye1sjwxPKGw
iH67zDTKdD+5OkM1z1x3MfSG2eKrj7Msl2ZCVveKrIT3qkXUu3GErr+XHluXZ8xH
H+Yb1NI5nQ+CF4aPeFymVAwV0PEi8LSxEkFiPW/x5OnYQg77Oys0xj1e7qrDF+XF
yAwkLGgi9SAKxBFiERdOcwPCtKNFWYg48aygsEs/G/Ltl+sKeFkNlXzy8gLnVwN5
phgEGXz/NbG/DOix5p52XMqNlzBjt+aPfEHQlooc5WZzL6WnFvcGYWSPaXCVpk1S
iL935PT3P0toOxYPT8jx44ZbfTWngNufEpseoJ+SjD3zV/qCTVP+3vW7PKpsthDI
PQ0/+JtjMYyC//4VdgIxUNe8KLtOSuEyupWsviKlPN40IIzIpnmnvD380e+gEaAO
XjxsRROJnDyDYyFYy6BSGH53D0UhLFhCgqSGtbpmByu/Xb8jPtcfbTvVxB+s4tNm
XkpatpZQI3uphdZgYfU2Vg1Si618fd2/2D7caXK0fJCwlRzWYAFlo/uBlSZ7kGgJ
v20zBETX+yj+dNz3/uEUrPTTtfGe6ZHOL9z0AxPeBGV0v3bHZadNjozt1WvxunF4
175RyCjzHUuOHI8cypWZmNOTuU601WTrne8TGaUe0QZttNdCZGFSgVCDAyjqzOs1
MF+1O7yVLwSSKM0Z8Uzgh9V4Tl0YQXl0bM4kK4rAVcypvVQN/LzciO93Obsx9Xvw
6bj2sSHRwN0JRfaRyX7ReL2lhK+sxAaZndIutTKobdrLQUOSEZUCw0iffJT4ecIs
KaBoKmOBTakcyishNUXyk0Ac5sdI/0aAKGO3haV47wTGR+fgCCbarddpwS8iz4G8
DrUBhWelbZkNR4Mj3Hq7xkhHtHykqmPzNEr7lV2XmtXNpCYoAIHNcuAaJPhIbMpt
VFGP51Ib+IYbFv6ZTzrEvy4E74fDBDU59RV4vw1lHNqB2GTaOevK8UyYo+si7VRA
taWiQ5HMmPZy5H4qi/XxkqZxxoUTkz1UboEykQgIKFgAktL7yG7jTUX+drM2Lzx0
ghy+RnPcyJlr88rKZEU4L7xHvyoGVvskFGR5LFY+13KiGDCa3Y86wQcYSOOyA1wy
rfa4wV6HjxS5o4ocEo7N8sscW/Dd1WnVedaqZeRwiiOuHl17Qpmj6MvX+lZo0Ugs
zgxP62GbtQcUfwTz51tss2pF58QoTvBx7LdlFTMedKBbNlmk9s4BSqU32MsDRRN0
MBkEgke3l9bIvozFonTYGqx8k4Szja0N4N2IGeKOQMG3aBrSgLOX8dYDB4wnfJsj
fjdg9N0oBMrxQKjWyDV0eXuaVklrWP0Vj0nRJvJwIQfYaYqSOhjOWPJopP24OlIJ
GL2ziW1Qr1NVr39jf8dWFJfKZi56UWotKdvrgin2MHGo5GhP8jmadZaF9wL+zdJ4
YORKzZYTGVGrASbYC1UAOIzBWAjdO1asDgMCWzdMTP5+MBb7Ht1a1dMXaksxOwrG
VpCYsyJRUw1S3b+fUv8/SarkC0rY6bJ1rK58xFOjJbmu8pb+CZFhe4Jn2KZjJD7W
5WNHU6TzIKFOWlmCvziMyCJ7qi1GKbp4CX2amV1lH49tENJ+ks4iHmp2r99olXGP
7aGSeEPzuFEf14H6jVicnfaq6NdOxN20x+3nmHYhzOJGigCDMU6dmVcLG0/HEyJB
VMWVCB67yqBBdAvYSIrYbL4GVVRmRajvjrmFkyJmfQuGAceTdtL1nI0Y8tVLbzER
Nik34ejYMj4+4xMHGD1omk8suGIuLIJUH56XlTqvjIYXO/WiWVo4km3fhqT6gbgc
A0rhtLZ7Bze+dXbRaKaa34/W5WHrDPQMdeCRy7oMKNBGb1tojSytTniNxz++37uO
us+C+07lfCC9HbMHf1ELvPCMwAQSB20SmeRD0WEgVv3kCdFnOwW2eGQ0X7iUgfR1
xUA8Z2exjNIYE9pesiQDSGeQ3ZOucjthf7JcCEBvBDuHPCbbZCFe9w4j8KL93uKF
KDJmTQOSFXlMQyT4y5VFIJi3g9sK/j/AgZgvGoX4gw0H1VYGwwW5syDsjB/0sd0h
rOGRd06DHIHovjuBvGPpOsNfz4pepeydftFtubEdqNBPME7rXg7/wejMq8seU9/A
o+nbtTZKR58Ogn7O5bZhM2PxU5yawsMpxQMronYn2PI3G8sYMaiTlu13E9oDoe4m
LETgwHuHC9npVsFCAA8qVRc1vQ+dAgoEZUEG2py0PnXSTvWkyFLpMTf1Geui9w4s
4FL92tP/D8mzxhDOyXN8Jren0bd5JepCkX+pEYs+9zrOaSAcg6eHM+GhOgtNFq1u
x1Zl6v1CJXSM/V7ENTH+d4ESMUMAAoYZ3vOSKJFxnSqMxJvJdij6My+9zB6u1WMM
3tTu+h9DYjTYLK1bFlfPNADoO/SNDGITQwBNzg5U7K5G+BMtwqhVwcL1Izf6wTrD
1zBqU5lPTCtWHmdhCRPBRLrXBsv35aa0P7gHRQKpvZBddYlSFzBMkNPaVemn2gc9
LWf4OP3/GcHpebjwcZ9sDav+2MgOS82qWC0XYNvgRFq4DzSd62U7ypyzomSDzUpl
68fjLH2ZGvmFilSo1Ef+5VUzZ/a7NlY/6yhgPyo21nGGWb3v8QmhH+djsAhS7DUT
lsiL5rAjZYDlb8pxJ8EcpjcW4n7bQtgGLbSmppU2Ypt8AzmJHOlKkrNA63lPIXpL
p3BptovH/ATi6+6YFr+SbbOWOkOlfECXbueOGHlbqlnmaw9SOYz717pccgsuYRwu
3ULysqgU6ygNpkm8L389zJ8vobW4gIWAmLbCkqF8F7tGHGoQxlmPqBBtN2wmjy/Z
5ezBRjbkpXysvNh769VRlzQV1QnVZsOH1WBJKIdAYRe4+dD+3phg6w/3esE4MkfL
eegFwKBhyUDEqRY6O7Xh0npb6NErlfb3D5FfJDID1NLQcxdqr/YxKLpCJFbonwGo
kPZyvdtbWt/OO971qdTf6IFSaIvyiE2qI4IQE74Zg08rub4k+2biIBb+/E2BhdJc
8P+wSjfJ3waVjCB6YxGdxBHTYSzMckiGRESMqFKUnFxTi3cctOSn3cfF8vgY2n/I
JJxWF1xUr094b+On8uB8xSpMrX6MzFXd67ojHPnMXuJ8g8PJBguSOo7x986e3Bbi
UgUaSF7F3K6R0XNYhBX/RSVbiErkDkDTuKAvSGEa8VLC7+Dj+vZhxbmvQC0b3hwH
7L6OsXJxd2cwjWwofcSbDvSCXTy/14nY86Nm/XahECvYizqXq7gqqUVwTc1s/6Z/
/qtf20Vc6szv0vS8UNZQ4UNAadA5fXO7VJcZih1P/rA0cORoT4CY8bdJIxBo4Ouk
CSLVs/51KxjMufU2bAmiYMeldd9oAb0SNEQW8IO/pDmsiwEEnXaXpnXIX9ATCG3T
gUZW/PHtDH2Q9E+J1zaa8ahOBm7wcATIktihI3Ksf4HQuk/F3f6V9DKnY88saeBb
ULln55MW7eQ+0FEEMNzxj8Bj1YzaRJqq0fivUGg8Sw+TM/0ddqIinAsYmyuZwu+s
bWt8b30Mh2ubzJs/BLQopLqsi2rHE2xGO2y19gxdch1IKxGNPf+q4oA2Abta5FuA
hin2MgDhWyDKLzdE1L89WfWaPHF2a80os6YDrL6onSgTbbxrKncS59URY/eYkgps
e33cLxlhTRNfwcn4dddnrx9AFGctdt4k7JChy2tUHUa84N1M5FXoV1LggFlV3SC7
1XTEXaRXu1JKvk/dyyhHzuixzYVgy/4k8GRpEw3JvDYE6dLLfRmv5YMYP9f0Q9HL
MBplv+aa1IsqAd7Xm6pdD5ILOq1aacCtELG7oRxfziU+6SPZ9yQvOtzczsjxyzTo
OXFf5DlkAqsvVBGO3Tt3Z7YjFR7QEzYgFPQSoXR5GNoA4uKhjt1B4faBx/4f8KUT
qcIE0zuWdXag0uDWZyzAmU+IKA0LR6LyBB4CZ6DpmJseJMRNuCLZ+kHb6Oucsmak
gMuRcey2Rt239lADFDUKQs6ZAkJK3lSHTdy0P08I4XLNule3SLPh7l5FXRtuF01t
MLoIHji3qC8Pb5W2KbwMb8tPIP3xYbWnjgP+NWqREGiaiV+rntXG+qEkbk2EWs53
JTiVMdWjvb6iPHi7Fw+yBMdZaHeR8vC4LsOSZxaXGUb94TkMsktCpJZbMGAywIdu
JeHrOg+nQSjNtfvGyX/R0yY6O02aKsAJcq0hGUtIWVHsIyQJrJxT9G7q8ecfk6Cq
VaVTfAhJbuaskTMcXc3b3W4EBNuHWfq+1D6gFBWNqQDS7JwRQZH5RPjnIkH5HRt0
0sFLlEvlybS/bBjlNSTIptdt/TKqxcip2Z9zyJg+Z+7vQesxweS/hOba6F0abiHm
Vzrp6AS0IM0vENJxarv8zHnMLjr0leAY62qksTEfS5qJSi1FmVHINDcd8iYIRmMS
nhpl6HYA2G9sagd4LZjWDQRPxN7NC5LDouWi0sG87md4gd7yFhcYHHl2tX1Nq4dr
Ic0y9JINSdMWCZbYDoaHs4tOcB4N5UjH5lSTW4MnU1UgzdRr4dnB50seIZtU9uBj
hi+mYsqzQ+Qc3F72uXaQItHaax52VDcywmYKerO/xSlbsT4BxS9i+3HdBuyXkVXB
BlzvEQcr6ckj9orspg6mvfXqMP/GQoVq/xIAZ280E+so8DmUpOp3T/oV9/BWkNve
frtFEM6aTdm59hT33S85uLHbdicX66vQ7+NzghCLz3CfpTFPI3q00zr7P7+6VNyy
K/1Duq/zWSzqTHGHZD0JLZ3aZsDEZJoJhYv6YFfoovIlPB61wFZSWSKPa41qwggA
RG6mlj4rCprC8wFJZIgMdRZKkRMq87BjInaBN+Sn+qOMjMAekqpN2dFcGVyDKWjm
pQGr3e/YYY/V4AY8UijZzUcayCNusR0hqViERwTH005q/Hlx+i3dCxHGsafbNLKx
9aUl0iBqnpktKConfc+kkqjd1FvBGD8li7ntxmGDUNcopkoJ/p16H57uH+wFwJPl
7cuCbs6dPGom5BtLrTmAw5eLneTkZgIg73nhQ6eHs1ppYCCVXAJG+548O0dg3QL5
fk6uj9Cu2yWKfQXnTcpxvjQfJHGtbNU/boUp+A1UKm4hINg0dW09hnxKRj9Pd5y3
gHiNWbVxX3wKDo+YZ4AaSr5aLJtUTmpw451lhl5l/ZU=
`pragma protect end_protected
