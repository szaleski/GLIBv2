// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:58 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
TZ9D3ajh0Ou9SBHKz3bO9o5Faf8Gl+RF+nmcMMGwBTDBhTw17Wu6p0uEXPJ0K8Sn
MseMMFz56N2n8nlmHh+PhMCKZnZ0FljFXnyYRkOdAWDTO3d1/Dkcs3uNaMHtiZrL
1xe5d0dg93Q4wyaHuGtLa6b3XnXFEBCKF5hRQ4jHjOc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 21424)
qQez4N4a8xmj5FQImS3odoX4yrP/D7piO7v3OcCqSYnVNUexiPXZbCis3dx+4pwi
Xte5MOoENjAfas39JqONEZ3x8haAUvJO9m17s81OX4An3kgL5x6VGPmZJH3ey2Hf
U7WONiWePQIRBPpsfMYu/PkCzQymys2+ioNSIFBus25Fhjaiz3gJ0OAkB4ZSo52Z
gfPA5TrRcy909XXzXnyVUaDaNpDaZdLiTvyCEsNiPYxbHgZe6y+flbSSOPRY/u5n
u+O2wvJli/dvHTenO9JP5KKOgpVz/aWET/ar14bhuCKGZ4uATps3+4h8yy78AFGP
B1NEhC9yPDFgeCxIRcS0GaJRUfeZuVTcr6zgjTm/QynEtqEx8YmBrFe8qjIytxHB
tR1nfhiXOSL5fhhClU1Tsiao9/qZuMYiXn8bFq8wY4qVa6BDXybO4Wf2TR2gEjx/
JCCQx+G9dLD6xseeDZp2qDvsCy4um4iEH3ZY6ec+/Eg+Se5/ba6LbjIc2L0vgEDm
ZLTJ7QTLS+uePR14S2DNV/7WZoCV4cpLz8XMk9thQRlH1zB4oh5iP3Un8PzpJEXa
UyKuGgaqVg88me6pZ+B+2IRRRIx4z1zlgqFtNpKh2zKMxESl2svYU8ppun3g9NPl
yHWqUreuhTHpeLfykc8o8Gs7qPXf4IZ6XPkPO9UY0yY9dGXSzppQelpK5HiIiu76
2kSjgdcnZhhWgCaVAjbh/U8OrxPSv7ZzhOshVzDJC1/vSzErX2vbYv3sL9vQTlUL
Xa0DY+v2EwJTIlgxzjLBjvWLQTp7jwA0MvXTWLKrAy0cS3kgK71T2RqvLf8w6cNn
v9RJDW6kLY/bMvlW7QzHWzWEv2vnjdyf6sLdCWisdQTUBu6SDk2e4k/g0NTn4pb/
VlLW0FWXQvCyiwtHS3xPsueZ0mmNdFwR3oY7KpNoWw8hTyJ+N3S4hAxsJCzLmyJ1
FdeoH+OZp91/Hyk30pGt/2CMtWD+ohCniRAgPPDOeCwTxalYEst+iAXFLTHcZdKF
xQW95AOZDx+SA/jtQegK3y7rUUQ2CQc3rdu7a1GSOTtZGTYilR/MyWEODvr/6vjQ
gg071sj584EAjzqmNdDPZFW33qmhke3Y3u380tnPjFJXyCeAj0nCa5daNigz7Y3x
9WhT91l//E/VKJZWa+FRK1W5XKpMhBmrOCPAkJrVDFv1+4rXPMyYVoU5i0x8DbVS
KCua4RpT/EEwPysKbE3iT+1jPGkcO6jJKme0biQEc+IXLzk2p4QsASBpPjiLe9+L
7RRcnq/QRBnl3QIs6uWc+wFcuMe9eZYUGxmBY5V9/OPMbKsM4BwhVQTEz28Dp8+3
3cevHdsNKQ426TjwIqjQlabUxyQpEYFQVkBKlTG3zpqQ72yg7go0usgAoSciwewW
Wyfg525luInJbwDq9uw0RUJ2XPOT8Pkx2FJLBK+zs1QcCxouKfiZ1+LnbaKTFOwg
GmSgep2b0lDFh9VSrTpSTsyR42Pp9iHQi8ZtCy0pnamrdDtKclroi0Ps8bKOzaS2
IJG3sChBoVVCRuJBW81hSUtzyfe/agqzoWNr9YV16P2gt8Ycj4x6Nc1inyMvv8Wg
aB+QA90zLeIzFI4X23pG1WQk2nStsQVq6uzLVy5zs8bWS7SNGnCRJFLHPseca4fB
IHBTHJ+COIr/ZfoO8HSq2v0dIE9sMrcnGtIgo7PAS6uj5A2o9eU6NAOSqjYXSKmm
6wGxU/Av0zJq2QdkGXpNfkGM+ZOfeaGjZTIZUgjq2XNBv/qW/JIzBFJ3ckcWZ/yN
bZ+NSPKC02NMaoUcw5/tueyjgwjSNZ9yAeyTnR2HH1j6J9mn61P/nOukrzroSpeG
sqkbFB5N7zXvCdRrwwZ2RwmcyY+p/mM6oHR9OTZwr3jXtJVQpFDoIGMIwaogt3cB
QIDKwA3v6m1LHcCZoA43yqO3Jm75xomDjWlHEbCE4tidNp4JQ0DO+24DRHcVuEgH
bvyDJZTDTFI3aaOcUNelguSh65eZgTA2WqJdI1ALVSeKQF+alRuaoFa7sNZNjYcN
oTye1KuK5TVEyUPFS2R03t3d61fGU1ykib0yBLOj+Dsx+2rOhtYkeVYc7njSn/5J
2GQ8e7C4cqVaFNgGjtp8mSDXJaW9FC4gl1WnRFjB53RrDz+bvTFDm+CZ+2HwJswJ
lnebT36K1jwOzQ8pxWVmHboBEM3P6qmb37L2rjSVWEdi60zhHhd+QLJzltc7mwEH
jvQW8Tleqvx2snMyBpNf8Km8aXp2io9V0YoTiw5BXGmZU34WSTlfBSwr6bKi1tKK
c8PwsbFiSxGv4/wBUiTaZNzrH4G0IGkwAf1sVZb6u2AErApY3rKErQuaICPn/Khk
eWxxGuXVFmZOPT3s4g2ZUYbEL5dUpq5dyk/l0wSTMpQ8w7BcHXbTJbJEpfKx6v2j
hGiM4MO30K2HD96N9s7fX71KBLbKixasWKEYNyON5tmXRBS2X1BuK5DKOQ7IGUtG
dWveDBkHCC8HUsLKzdrS+EGgeV/396Bd67Ra9FGUA6E5UsZD3et9aJd7GGBrpxdt
lHKOHElrIHzjMNj3rIsah9VOnrzdETPDabm3ppkoFCDvgN8q7kigyaySmSyVvA9U
2RVJb2Tako8atnMUNJHkQOpSPVpOvS84642LHTLNPvuXQQvpLFSTXZSVbW94Ir02
YUmxKXtznrR61VDXItCITytKOManSgHYnSCx+bsrnqn1B7s6iazv6S6iy1++tlRU
1idUhm97hMmCGkKSjJxciyxPLuZ1lUOehhIrFZknIQjBIdsJSFNv/Z6DG8IhnMqk
3Nwt0JhPxHUusi9HD+NjRJ27Uk3A5De61ROsRi1OGLaAmnOXqiq7dqZ25rKLvti2
oBkeY2z/UgNIZ4NMYGpONzsZC8eCXKhHz0MO7v2JyqWld31rL/eOo5/XOgLGh6e6
GVnGYWJXbiPIGXc2u1I+fRyvwoRANRmVG0xeHpn8i0dSxTJiwW5YPa5H9EOmi0Pa
E5aXn+Y8w1brZM4OiGE8FYfLALYfooEeS3IznbnSgJabVb2YdTES5GyElG51tkYn
u/NLHQWI+dXp9RDzRn2klRMqyBixwv8WWOc7N3004zYwVHncCjEsEIQOlUz+7U8i
qo0aJiZjnvqZuKkLEfsAv9ECfpcE3dDH6CdNNOYUDXU7cgSVVoM8VOtmMYzuMqUh
Bs6Lyuni24j3rm1PJX6KtTGswDh7ma6wh5kNYvGGgpljDh9fGmcYUyIDXQX7I7ju
NuBEvBdnrC5YyV28wRmM7vpeg2gxqzz6oB2MhvGXIWzk5sdTwLdI9f08sjE7XoZm
9toCHmDuxhX7c7xN0W5MaTxXLyb7DP9aH6mVEbx1YidMw+bhHFLbsfgMoqLPwIvm
avpF7lDtadig9R1ZnDl5o0MjG9EBFRchV9XK17i2qyYOwBuVptiqc86maj06LodQ
UYddvPDEkcAlEIl3Z08Jb4c0qupoupUqkWCIEgjqWm917sqaNlzaE9vTfZatPcBC
BnOc9/T8nLc9c73e7W6ek2GnoP+yxsYY9FLAbcis3cb8IDr0xwQ+7lryzhAlVQN4
9KoflUCo+p3b2EEzScWAFY/PeCA4eTfmrrAvkwTEXhS+ZEz/xdkxjpqPCpGJvNLH
yBkZVH0NDqLQsYMInl05EWPqSMpWg3Yrgb1J91BJKevwvTfzF/x6LAZ0c/WA7BaZ
8Jx29UprZMmz8YotNQPI2ShEpEwaKcAT5vmtypwtaGom9t+VCxubddF37/88jMpH
PepJbZ5AwZkHp3C4DVMJY85ILBUpipmfLpAD2olK+GKmaFNr8ST2xcnp0/6/Ae2U
o5VZ5jkuozOtb1iscT6nTmuLwe2aHZXu2eDSHXejCXJl1krowRaQdGYYXWE+hiCA
B5Dme2gD+nmXbHgD6RNMBAFvv3QLnADxEOmeClUk6h+HJMfg9wcSza2fWHFkWpB1
Li91hkgw+nHtT7S+8iDz4DaHvwAnl1u+F3DHm5XYivloWzjtc9I5dFbn1U5wMHb+
0YOFww2POwS1mtX+MmclMXKcRG6GqJ+o+MeSLH7ryeS9llZYX7pvq944bvbJNrOa
Cp1j6gt63wKlFWp74luV0GdyCgVR4+5dUsf4m5932q0oQ3mEYMZHRLPPWazdTR9b
kfKRm0m3Nk53COxIEoEbNWTfw9LDz3kl/Akcl6nHdG1QT1N5rLfr9abTs9bpiTKL
n1geN/F9AZGYEJ6/nXta/wh3phyWHB/1s+LPrGIHkGgR6mn/GDwPkEKXiT5lpyTx
Ahe4PLXIbMWyeFYFgr4gVnkClbhuDM+KRJalTVHRqwNwMtRw+hthqerAwkvD1/iW
eq0HrW2YsCZS3S/qIV04SunXILaf2wveGPT5CYCx/VvRHoYNKaw3mgLCSGrQMJ6N
xB6Ax3hbAh+JmFe54pajydLBPpJUZvTWo9grVK3ij41G9JJriO49cQWaRQxxhxqn
8cyLZ4NSHD3atbs/yI7/P9B10KsRCFUfv6O5x1CuBqYHjAjRI9xIkfuXcYaQY5VE
q/qnZOfg8jg4Bt8KaZZXsYyCEc3HsnoL5MbMHUpK86FrYv0XKOcb9+lLTPkBCtny
0s0x09fF8p+eg9WU/lzBPw2l6MebLBXmoEmcCN+G+OXrluKHASb/zlsrrqaZStBN
kjVZho/6ZnyyyRgxO3/nYxRkccniWiVHdjpbYOgEyfPGY93441qOMbwc4Vu8xGor
9h65meGpXNbjRRMEa1UJ4C0c3bpoBiWvkbqel9o2J02sGCEzUjpk2n3FxLQht2do
tA/+OX6dnH4CzPuPno+xkVJeU0zCcCetdT2+s9ThNgpvhFOG7KuqVgm2tMZZ7EHX
W+4plV+9bMrtCtXcz7WZ7I1bbwleVF/PP476d4N07mnLslMzaviKJYW0qFHrqRBf
lPfulM5b3qLsr6O19yVKskfwiKFqTRAq6ahLOKI1QTmxGqcfVvlL5tMZPiev9/F5
vNCXHiMSPQTvtpodTHDgk53OSVQxGcBVaYtAXdKNX8uNkoaAyifi3jQOVaE8Wz1v
SnWRfMrVISE/KOiqbBI4rwq/MtTKPX4v3EjUhZHg+9S0rXjuDkJgWd95zUbc6hAR
OSlchzEPUaHIL7yqT/z/LRYMmGcOnTPwXF3XEcx5bqeUOsbiORPFPHxpe5jaKcGi
5kyW8JohQbDY7SRrHMUQWWUJ4jk3E2MnuF6YbvUyzYzZPcmFaxGSfBjTAfMlQlXf
XP9LOHzRri1Z48MUQyokB3NOmPOzUVEhXKY1qfCMGL/S4a+KgdSJsRLBypDG9U4+
aczs9Hn1RFLO5vnMPMRFOdyFOMDoy2FDRw+NXcEhN0shdAA4kLTPoLx6wRfRvQpo
rLAeyJv/tIFKASywx6jBsG2FYYiArcB+65UxdzDf2wl4YNvJB46n7VQls90hQ4aX
svCUUqJ9Zds/hdG+dxgSndUMjtI0PsRFB7DWAZ6l0kn6MQCLxDKApsNrq4LPSUGL
kqCgppog4oLrf6I9906vZKOk/vQDENhuWaJ1bjbKkkZ/gT1sM9nY1DtDWaRKyeZG
PuQeSW5fb8+q2l4N1/t75K9xQdO/wmTxJ8MBm8Dpi+nVCk3/CpDt5SlcQe2HY8j9
CTeJSkzWt1YXNhvUmQCZU8vBzFP7ryfz+4ZX7sg0M+j85ceRNy/Tnk4wY7DoNI6C
60JFdNHwuE+4wzPiNsf4AgpyiP2cg8JGy3ggFi0VLqQ+YHs2Ooo1T2aUD7OLom0w
Epo5BBp+LOg7gq8ZTb380PUF2Kecu+2s+7wBf4EJF81mSW3Niaj+nWGDej0K1j41
F2f8v1u9WbdvptD5gOyvlJxAzmbNV/fRnl6+AO3HaRWFGbSY6q9TKZV1XvwDvPFq
mtSL3ggWWUFVjDyCm4OmLb60ZyMytrfRLRBDBwgyFjl1BRwcrC+bRIAml+/NsNVG
H1fIgG7yGmAPs/GrY7Q9ZRVoEXHYf+Wpj7yrBLQyymr4lzwqxP051xWHo+ApTrWx
6KCOrkHdxS2ei+UZkIcbRdd8CpCx7aiv4bw7rCHtim+cZPavofUO20Yhc8RRXz/F
aVM+Fa1h9aRfqLBAEhRRp35trRiGzLeg3QO2pmlWsjGgURuli38L2i+Q0s7Ffanr
fJW/wJG1jTTo58XFgQsOXqVD+CsI1eKD8mUlQivTybJ1IDt9VAic3v+6ybH7b39S
bQtofDrEh/dy6wAqSx6QdkelIqdOIe705c3cn1IBElh6+qtrS1GkHWIn/85zQSUr
oRLoqszGq4X6qBwwbN8oF6oKbMuZYBuHcyvxs86w5veng33awR/PIF30wMi612II
CEkWiLJxORq46DTF5rs+BO6TJKadlaPX3QYxtLUPYtAPW1Bk4JXUgipSzblkRTLn
yGgQId2/AtXZ1sxDbr1/k5IWAaXt30Vb1LuZIAiWlsb0ZCljKWfPGI3AbM9jL10w
Ba+S4pSXQujr+ylctx9REHFsXJi4agL2C+AmwCi9It33lWvTMMhszL28N+U8qZz6
wB2e0Dl9Me0XDLryNOOG4NA0vHyMLRvVlFxa3eYzN7EyULO6QPI8BqjLMLTwl1MH
gKD4BZ/SUGIRhUBvy2w4A6w0T5W6CVI2ofhdZnZoMpVDTC+3qwXPknAbzf3Ne7lP
evcVfsPovi8yosQS9xa1KMFnm5wx6Bdm3Dbmr+6Z9l+VrhDssETYQOieHq4FC6gb
ES1DTOMd/pmbrq9eeG8akFkD/AEBqL++T5VHcA946lHlGobIb9XcNWIuj1ypErPL
B0q6lZrFadX+Nx1jt4cmdpYQWgrry+YzdSDJo7qCigx7WGs1vDST+EMhhnNbg2gL
V/OsrxqBGza8ZVcfn82XoaD23E+Dqqs2FdYkP75dMrvHSEmEabNHMBBLi201tx3s
uNY0N6eQ+2S6cdhuajPjCV9XQnEHE07f3dgGxWvI3xWGhUUCgkhh4RE1Lj1LgJak
JnLvOE41BCF9h2OJAc6Tq+1PE9+m/dY7sYAUwMOjw97gblW+b+nSveyDJGck4ukJ
5CGVWULsBu85LzAaX/whCpA3La3hWnDdeIT8wfIW9bzPrl78CQQakH4UcXmtJLsg
TB1s7dDWeFa7Jse+iBtMgr90FXyi24eoHfizQw69XPTBsj84KlvQzZzm95qMKjmm
WhmdsmpUBo0ZtAKNW8s7w+pwMTjTmxc/jwyS18oS1sBqDk3hieKSanPi+FZ9NeOX
P5+Vd6XtEuajl2RliDAHOaJUnXj2H0T8yTSK4epbyGk+RaHMUdowc3DkpdoD1ilB
seGUIS0aHZZNwnKSebKbuxPSBwRyclnpRD1QnITMono8ZErXGrsCiI2/O4UZ7fsl
1/yFIXtNUkhyaPd+LRKO6YIboi9VoRLQimrtUit26YlCgc+B9nILcd8igRxUxBQR
HIQub9jXL03wPZyO1BK/bTR+hhRpZ9/ppYzlp8f+wjmQRvAV4RKdv+keSRVF2Iw2
I72puhRUGhEXd9rbw56h7/Pk+5rIAAh1dOK5EKCYGhUndrb4l0s5tui/8CdiOR6A
hJDIY+sfGCEUXIy/p/FMBuhbIz6UmzXmbOSkAXhUqfadVBtqkiS4xp4BAB/CWT4a
qqnp6++mWmACp83Yr4NLEkwX+9jLpfNbvjGzksop2SXmisrlzzMLfAHsUlI3N7XS
AreGZnxj6l3bUh7RbL3YZjQZQDFON1Ca2reputfaJXKmBS0VbgR+ZNy2rMUiHGEj
C/E339Q+oY9hffv1DyJ5k4ANAg9CLgsCuFJNM/jMfohktq1NtjQiQMQ7w7zx5wCH
l6bOrZFAYJlBSNCBY8DVn9Yf3iFsOv3OGzFOdnIHMeAXmciSC/SHr6L2RHdPIAVu
r81K5e/wY9BnqM21VrM+xP/IAn7FNWEQMq3mG7b5T5gzHZ4efylelmM1Od7KlT4K
S66jBq09eORUTVAIJCmixX7q8B7CXrtD2h947OONhANZ9AhEaf4BEzKyuzUubmh7
HtFYFiWjbJ8/RNDN39RMNJoG4NX+k9sAEahiFjqKZNjBS9mTT4GMfFiV+vmKG9Dp
XsKeNqx6eGVGrAcz+MxEynSbsIdK/5nvUEG8YSk+31ozKhIrsad58C67NHFMad8y
tIAI1i9kfrWKnYBmUYn4HW7YUHAmPx72AyK3+pclEw/tRUaCvxWgbdukY1HATpEA
UnTbQ5nCakYsyRrjKSzyTAMSakTLiM5m19g4cB/jYEWdM0gj+cCETo29tRSEWMHU
+Fd3XwFQuv9qbQuPFO0oxTQQoRU4ZMAltLXhps3yG5WkFA6DgvRe5Vu88J+bmg+v
ysLXodiX6PQSm12uXU57Swg0G99CBBWPur0zQrz+pacCXV3Lo9j4jGYxYGgPus74
0O5TSPPV3IoXApTirT8RlL5oBKccfSn7pUGvkhJRHy78Kf4Z44gQAJXW7ESVmSfy
iEJk28jsLbBKr+JvGHM0UFHkaN+ECivqj9zTcdE9vFG0akz93k9UfRbjfoFtki62
DCNqfXBpfX7fW1rhGUIVKFxsLUwAzB7y3d6aLqcf6SeMY3VGpdf25LFgWcUIdl2s
+qSjdjJPyoCOWw5Tdbw+6y8uiWTaXN1mKfFGWUozedM/iZi9xi5JYAlmZ679kAGU
ven/0PUcb/S0Qw4A1+feqYAt4Fzjtr2Ndk+ufsW66rjJ9WeMZhj+r0rihY+m/zP+
XvyCSODJIveTSJtxrSNkPWVlEyZw/Z7VES8RT66ML3LwbLz7KMquznwkeKMaDqO2
uY+RMTs5UHqUn+QpNbWXMjUpcz2DHXyzCCIN3pHyahdcQ+Qbh6PiTHzATlwBrFGS
8gunEeY75M0ZlC4WiMJBui8I+VhzbfUmq/Ws/td5YJAOYTkSW7WRqiVCAs+MO6fr
xKKpRbFBw5Z6CeYbXhk13iBGmHgE/mXVskLZCJe8aeOc0Pm2cXafR2+4ReGIPbvJ
0wfIHQ7KCKTwS4xCI009WJiRDeeTFHB7k1w25wAiwNczY0eBnXQtWXqpVOymPqBf
olTi/Y+kff0yVcIzkDOCAH/KqtZf00bHsuMrlL25wClEIc38SOiePMAjSbwsh3j0
MRJD+94wpWJ3db3cOzR/W9pbmUbFJSART2NuAi01zlla4k8hE8iUHN7tjhpI1H1M
x9gpc9FoTCqnfZFGixgEWiom5W7XoJpo/gcbINHwELxyWgyU6yMf46e7ngrF5Yyw
lQeVKbJzaS8nc/6ENFsgrwcVc4JoXVF7elTa5NtlT3j476i1UNgNG8PAcPC9GRHR
D6jMngIgaHSEFhAzpzD5pjWJSZ4Xrt6+r3njwaxo+qViuZLWEpgIV/3Y65hn4b2k
7+DPuEJN9QUKTTN6D8nV9ZuAFKpygxspaRBeZgvsEKU6SZHInFjdsl45YlnqV8t+
QvTt8kwhYyKQMsApasMrw864nHnjylq4mBUz/8e0xwcZBa3aHFdhi6O2fZJXkSBr
uVUdXb98yuOEjUgKovlW4fw1jCWK+Y+hiWGyV9GvkrU0e8SRBJ0n2mBDuT4aA6W5
yiFgOB/aVkdIuxfisuMyZAqE4MLeDJK54AWgLqoFpukYCxeTkOxWsA/BPWf35t2C
3+NK9PPG8D28qMDsmEEzRVCFFiBsJVGqwWJmgU/F84TqkqmA7JDCMTGDI/FE23W6
B4HD11aBO6chI9aOYhzyfWDnMPI4OmFnIkJOXnYD6SNrHJHUCISKZ0bqnihm44bl
tGCwiJxRiSysQiiSPULx4qQaSgFS0OOOId8r54dJsUs8kqjkokuP258iwL6jSzP5
XAZnzXd/aQkfAKK72c31xiaQU0pGjEjQ/W7P5HI0vPss0FXfBl5PYH8Z6lbaHy19
c4NVaGDwRyQ88QkoKBj5Pv/E64G68hW+pi84NO6GXWN8Y+KE7GZ7kD2vI4WxA72t
CmzhXfjObSE/ftaf2lPAo5t4OA5knH82kMTo/9Z0d0RkA+iJUcsJQAcCo7BwwHbT
nWMn78pR03AeMVSvRsCmBIB+ZOzec6nc1bUFo0JqDN+ghv+yMze6pIlHxXKCYPqq
LgvY6Y2gj0XgcP3iiLItBbhafPBNyw9FDBT0fc5Odw2KQYsrdemtfcwGgevl55WS
6pPMM8GZMtOFjcoUy9VWFiv3LZwPG3LYtv7OMvaC2easj4D6uVUxEl995veekMtZ
XX6bTBmcxnmdhVDM+o/qrylgAr9aGg3N0TYH+ni+C6swFE4FV4v3N2RCMjshrW62
MBZSzAF5C+nNZBkR8THpSA5Ll3NCRpc0drkJG3Op7wCp8fHeqsN17ceSCAinBHMh
QZW4NL3cnoDogtIbIcQzD9JNUhFyvElHZAPSLQpkzN1mhHvyE7eYwJIMS6hlz25L
0gTawhrLblxdfoR4dnWZTU7sKD8qC8f0V9p4/vreE3zzDdFJ0quGx8qLPicxeM9i
Nzh/TmncOh1Nc26BjY4+UFEmB7KIzAQYzI3ONwH6XV3bGEK73tR+GtaDns036yfh
yxYLaJLsEZY52N9YKzNYEl1VcOzMqF728PeX83ZDXIlwIcX0cBWS9rzOh/KOTrUL
RiHpoMY7HoKx6eEPPl3p0FshJka8kCJfqJx0UoHTiHgrA+N78YMyILtnx3A4C1Hf
j2fhPhX8KhcZ0XDV+XOLukVBQdnkXYMrQZuQkF9QtcArtaGYUG0qDM9M+xiczVXK
begUjvdttdg88QvzyCnoYAgV6DVVUvYoua4egWJ04o6yRhDloeNEtM5y3g6vq7YU
UXvAJSZHO5g6imAxCtkSuid4qrCZC6I4w1GKLIBGkn4dTHqmsmpJg6NRicuN0fkI
7gNm/I4gtcEJ3C4fxr7JHQ1NveWx4STWjCTgkQQYcI019k81PrrNidsxtmuxCGvs
2txscRUaGKrTJTg8qHBF1/AICUrm6a7DpoJz4pF2p7V1k1gg3WlQq5GGxavvE3Jt
B0c1iqMe/dS5ZnfVCpaZWGY7zOcNkKgRaDXv6jU/EjkV1FuUzFHAzwzEbjH77MGh
2khNXYmESzUTv19mtZTRCqwPtMPguDmPmtM4MiZqvcaSPniEVpzuJwRsJdPy0AyE
SuUtvAtECnGBqtwN50Xs92rS9zvP5p/bb2//OeR7pMgKuZgeTGmDCsWcddVbVyxL
fWb7b9pxMd/j2Ii4qhAM34JGPLgTVquMWjzO3s8ojorvZIscO1n93ceQiIi74g35
pEuIkkW3E0muyi7hTGe7jFNJW6R+YTbwXfURmVFUk/wdKxz0rGHbOj+cWiy+AMUN
R9y/7dsN0L8bUk0cWDAEuyfcX0rxzlMc/ZkCBjZrOLkLkqt/XhcSHPdz9A1mVAem
BZ2iYJvx80AKwAYtrfi3KYRtzXQGJD6OwBMe8cC75d2N/B9LUY/fUpSIsICWeWbp
vOJTIn0V2d/8sRwuwMHjz+NCrfGUmyWPumEBLLXYsjc5CA3scpMPz18pgN4/4wd8
cDaBCUcTm9IvoxCb4+Tj/qTqTnwNwGHibzduSI7OmzwLfrc9mAJ5IhlHb6Ets1ja
cXJTKby2b2RDlMj/fF3reOi4pOeKzunHcHA8XrZrXThiZLGCb21cSkV+TNrOkTrN
cviRifyjuSXL4YRk/1+9bO6aBIm5EDjYQPbQMbXWfl+ZccEfjGqALB+ojkriRqYs
faMD4JJemKItCo0twIRaIVLn2XhEK4jnLYLpoMsD3u81lS4ko0y0DgF6TcI9vxGg
NgRwiP0RTpNLkVYwFnBtHNOo4jQKG9eKul1MWwJgBXX6paCHZFRVnaxDjtGhJQEi
1NNy4SjWxYngPJyP5Qm6+U0p+UY/F2Bbqnl7t2u2Lm8QZDFUC+MsOOgoEqK5GJZo
VccQjgTTGL9r1Vdc80ML1chmmQK/ab5NdEbPMbpLXpO7x8UCzM1pkfGHYxmlkO6D
NihltQ46GhLvFMYAACa4ESlfaB77vt/6a/9zdoY0THyQUYB6fcTyJyCefVcbsgIb
nc2QOBJXTtMzPxPC43uM+D3HrTYqLW9hs3HTKMSsCTAYUN+pm8oRdNQ5xHoHgR+5
SPvR9jZ6Vxpkn6hqRjeA0At6B2s2K2/61nstKzTHp4gP5/eA+SByWhq9yB18fusT
g/Bf4yihPmNq4h3uI2kIi6E/BdoOlE9HS6PRFqEaA+EfvH1OlqSKEf3/rwPeVxUT
7AM/kF4nkYcYdJDXBQL22PbDHOv76uUCshmO11e2Z/QDPdts3GUis8E9GvpBhh7s
eAnA8ZLT8YYHHxVPEVMF9jRBxPKpxnmoXnj+qSdsH17poAfUVVYDbkTs2Pls0XZ1
ijRd2meKvtwjhOTGpdsH2jQRUt4EDcaSdt/X3FX/FoI6eC/YKPd3qNtHJ2FGOQvY
51Tj3APet38O9UacqEi5ECQGYsJHz/1GcyWUcwzSON7Iw5XFdISDWpVsUF0zZWk0
eRwTUCd2OanWY7kOcR6mWWYQ71VjZL9Bh2AbCfBIk35ifr0/pPfzpU86M24LUYfN
vjsi6Pd8WdgXS28pPDNQCdsg53Ka1HXCQPFQlfxEUGmfNGIZohng+JbeNxuMIL8C
VHZBnWn1+H4gV9aGPD63vQR1bmwdRXMn+DXxKRd4ySTCcYF4174ZIVlFRWWPPCc3
C+qAdv82dUhG4jD1POPEYwiDRhC0UKrDD+/nWeI9GUctSH44EI3ztSYxsD0BGLa7
AHRT8od9KyBh3nKeMmrxASsbAWbAivb29A9nBKVnBlagdU6VMkWDHRvt9j7rQXgX
bHdJTtiyvobghph5PifNZGVd3PFVrBIeV2aGyf+XIm/UOVtxAsUxcryWIL23vnNb
93A97jOApelvSSQqxKLgWLyOs1A+0+QUqJHhEP1p7RdejFaactxQs6nhcTU0HTHq
If9HGeOg3sx+MdFl7LwKDhqq4J6WMb+u3TCjq1lO4K5sU0EoaaK3zSNP+25FkKcA
hGLiIVjQGiJFOCet9mNBLcJzyEedRrb5K92R66ZFacyZ2rAkxnhViFG8mXPuzlrT
qr9k3tE+Z0OGl8+F4qCxQWwsxLGhYJCG1HWlJaDShoEXLQzrzIMgf7w79ZZTnPLD
U/QmzHzqOo8Y4NrzwPdpgkYtPyJxsDH8y7ZGT2p0tGQaUiIDoy8YrHuHFckxzScg
+VN22JYo8uUGPkvYCmQXdnbzOOtMd0orZcALQO4Eq8Q/s93GLOa238F7wg0dSWTz
MSYFNP/6+hnVHu7FIWHC64w34yC2uvl76Dn2HukSdWMTG/xZv0a6/tq3F8shGWgp
qQzRInhn+Wib3xtMYuEFpUKbnPBRJuhAKpmwQaNXPzJm7GH1NDllCRR9R/ff7G26
/hjyeQw4UphWIZR8J16TivYG1xyfSxKvM0oI6BY03e44eYbmycQTeAMbCH9bzCNi
6GtrQbZOfoTu6jKafbnkjyXQ32JkwNzw2J5G5udgAL1xDpa7s1T3uWhU0IrcXrX8
L0f4x+NXXnTZRIw0BC+BbrGV7zuajI3+5Qb7DvvJbUOaraJebEbaYF6lRCbmPr+H
KqaPhQvNgJUm9F07ydkb8+d1TyNeICxTFxpdWytU90jxZdz6kZHQlZLJIHzmPRTz
YFDwi6s/k6V5YUEnXjYoTdkqjMhCB4sGRgP4l4KV+xluBQtZCBqKlTedT2HW0MMp
9WQGBhIrwD62Qv+bwyHIytNfrUQN11G/abyFEkRCxwVlqefHcbo1f1Mo+Ej8oiwx
YUDCrFxI0zMKVS8/3qVXKVks5aqsTnc1OWRBBVCmbj0vvA9jP6O9ifrJ3WfQmFYH
qaNEz2eAnxT8cQyvoEJACt7QW9olirDorf9lRsTJGtKRLBW4Oc+SD6WpkVakBGB0
4jiX75xRwehRB6wL8ODb8khELD3hQ4SSXtQ4J7hBmsJq2ZT3iYzmSrwNUi/jBPp5
PfScFRBUmvAm0tB4ZzCmwEstLnQ6i6QcchXg8xwOKHwxEh4ZTWAuOLBtg/K4UClD
o7NNc0S4A0wmUGecVwXj+xDV27/oCwlhUyQEGur9F9o+RLcCSpoBpfnkbFDP0Jn8
MXycqwF7s91/f4Ub2yMwXy3McWQd0AXdEqnlLhZubYj6rXQ9SQTBcDPfkEfIKcZ/
3hEV0177pNlHt2vTzpDjbAHRxhPB2OFimUIKP7On7Hgv0e+lE44NjhUYv6o+cW3W
qmDL0kEgOERH3x4ctUrmqJBYfAnkKwBYH0TRCO/V7QDUJJAs2ukQp0lhqENGIuPB
qoCouWtCUAQE6zj/8Y3Qcg+kOOpv/LkFD49rDunM0Ql6VSl1Ry5zKJzikn6R1bCU
iL8DrvPb1++tW5LABEkBAHAEl+9EpSC3sXh5sF4hV7RRCt8B+Jm6mtqTGXFNZ0l2
JV0fyYa2uxeyK7tLUw0K8FhkBneEpTdkYxBWuPitdLXTewDNrEbFe96YVlR0z72b
CPfbXyjO+8YuPf8u76LrpDASgGwfZiehxpvciyC+bkHUhVcqcNQzSGVmJ0sSeDc2
F7SUe6HPXqYxFfXDFcsi/6yaIllVjQRd3EH2VngIbxwFEEStL5on9EqeBprAq1Hf
uyiAmVUcdgfX5+Lz/kXBAmv5XaM+S0k7+1eXRqNX3jAI8A2c/fNwcHwe4ojT24Mq
hiIuDsg9S53ZbRcD49E3UGVIWTUOoXJqZN/DVequVeIrbHQIUdBjIkjXjZMo4nsf
0eg5use0vc4ZADCIftyX2w/e1zo3saGR8y9HjDVIeu1KYBzpnOawVczCrxXXjWTT
Lov2X4cwxMSanfIrhxGPn21vcWxQfyvGrR9nwuYgTf8fgFPN4eHexs90KdK0ra6m
u5RjHtJgWjBYIq/c/nvIWF6xYjuk7I5uZayaGfY6TvwleB6zaEd67Q28vlKyUI0W
Kc7HgDlKeEsYxBJrLUEuP0JQX/WFbylpxv14dFAvoJbufOtm0iSQtpSPaAX6ZHCa
Kv3hlUqRUyvOEI5iDz5dA7ZY9Oimcn/7Zy82foheL/I/Tc6ibpniRlwWumuKp25j
4iBfsRdAd/Q760FnkJwJmJglNuhtVuubeRBfavYOwCrWt4KL3FnTCKra6npFQCpi
KSx4tlEjr4EVmSl4xW+1AaPZdwR/fXWLNrHeHEWDR9+af5t3B0dn64nl97tNxHaV
3MI5rPwea8fFyOP2UfvXqhnTvdu3hTOjikw5w+iCP7AFcE0iEid0j+iXR4cUkS+E
4T7pnhuwVkmAf+n0l5JzQrRIYw/8S+Si+7y/jsY8Mroip+ndNRNSk/jd99WMXu1X
N1FJJUUIh4OWaG61oIbd032D5g8OPn5zwB+HfqyjnWmffbg6/OYUaFjF2IgOeWBC
k8i1eG/aCBCUyCpct4dJ5X28IDrzeWoszCjhp2bYsXJSfVgfN7VnB9ke1CZmQc4X
TcsYvAMnd7jUqj1iNsRCcv0Azki0lYqESCR4ZPySSPuY7DVSbfo2WhZ5/XUfVKGh
QfTjqhXLTMoLdvp6GbC1VgVC1taY3w089rcLpMZoixZPp3a8qBJLb1qkn0DYq7Qs
CQNOCv3FiRVD83vvBeswog/rSyzSlM2qb9fR3LZMYWr7ICTddbHXbmGOBwofCuHa
jk/IlKY1Y5nOhhHj5knIx9rxnekBSDo9A06ZZzic3Sia6Xff08Tc1iR6QBV7vCm+
OvRhkmS2v6bEZkeTSgd/bh7ICrsgKv7ndo/7VP86hBTjdgIJ53NLnHhdh9XJWxBa
f9XBrZ2pXKyJgVdqdKKWsUZduAybj3Muw+31uMomqMCiSCMrGOjFaOG39s1ZMRMW
mArTiU1C9AppI3ubLLPHizKOHWt+TYuo9vHMkz/+pUA6+oILuPCH0bUgLdEqMOZ7
78HlPGEvowoKAao50c2lWYlKzr5K2XQ71XcwOKHloUjkveu+tpzoAMlGot30F7jv
uG1v1qZ5xf23ZywkVJAWwOp+24rYQufjbiUwulRsyAtqMbFAvKCRvsN1BliXWXVw
mOa9foa9yrF+sQ5jXN73mBV67eyW/1KanqDSRa7z5TNCi3ng+d/3wnaEOyF4bcd8
NRc7yAAMRjlapVzWJ/TECLHy50LfWy2Yth45/GpjmVgMqVarFpyHWTsvvBrPtuUK
zQVl2e/LiujUD9yrih8b12YfaqfBaPEByd90xJvDhibsNqfTz6w0Bz1Qcds4D1Sa
KZvF69V2NyManjyLKJUT/Z3IixIUjhYl74aOXe8x+2UCdncjQV3HrzqP9aOjNTTO
AVOdn9feMZeOOQrk/Ee0AFqNYodsdUR8D3Uiy8pN6rkmgdbW9OfT5uwi3SJRV5QT
pabzJvfuQdrXo/KMrfz0RRSrbEUIciIqZAaexwqNQwpskGkHKOomlkkm7mrTfVWG
pr3LVtppWWXG88JALkFNCFstPPuqFGNfYg92rsqkOctrE9tw6jRM2jEwPggRRQTn
YyJ7G++NvUkuRShpr6h+G4DeFboYmX5DBbqQa737opa4bphxJg1Icv2VFV6LnoPO
JhlHSHH/aACndwMzXpc3rVN8itk5a9qGvYYnZ7YJdDdYs/MZwqvz3pGM8l5/kb+x
8hf+DDyzGigIpCqzJ+C5rUvvomMX2XD0Ujl22MbYuZCEGR5vkbbCk2urKnagyDS+
LWk6lhvxf1a2/IiuOXHcJYz3TAKO7k/VYEXfjbHygLj3gKNYaKw35sTal3uTSvSV
NFg1x/S2dNXDXf/6eJ6kjm2I+onW2Mhut4gHcsPfVzsdtdsxMnqn7OC0RqwjTb+C
8fJcinIkdRQ03NiMLl93tZtj0EFYeAZl95gMQBvU5Zc1GpiIinRO5qnTBKKlwyg9
1SeOL2cDeivp0M/aK/RUbrunSZ4TgKpiRKhhNmH4jvbmaP+eb1YzNR/GonBo7uXK
8PcOEfpGtmXmAbT12rZFFfhAJ58fYF7+y2b3MBFQZyFDgkUGV98AgIQHbZsNQJ0h
0l2kOHvL7DskbEQsiBaFcoigIY0Sb5vMv0s52s/YHmMJ5GkmUEu32pLMWy0OtH8i
y7x8U6lQ+phZbqFlEkR7134w7jykUjtudOUu3xINMn26oAkOqebAsNS2gp1m93um
j6e7/Q4dVq2boFf76PgIKdlwCiZjtTpYxCwcxm4xekJfs/Amh8R9gIYH1Vs9LFm+
0sS5V1pqZZKJv3KfSPUpNdRDJH6XOwdvgAPWBpRVSmfk8aF1GUI9UIX1Njt+ESn3
G6TaM8TpN0WyCYMK7C5/bocgj65r9aQvFCbH5SO4SX/4kwQoPxPcLEZp3P39fkPP
KH68TUkpdhWJBwtZYYg3WZMj6Z3Qa/WcbAVUqcTWsnG+es3+voKza+3wmO7ZXdr3
XS1te9rA4oQ2OcE7xVDGy3wUS3o7UjKwEd3Pq9qi248kF3O0ZbPH8ZzPJLCTZgCz
lbfvt0lFeueKXnciZBequ4OSqIJ1wnc4tcBXehPPaSkBVP8iZC2rT41CRBg8PJiw
pxY7t7yehwzlRoeg6s+u2k8PIRW6MpIHlTnyHCZvw0un9v1PpBDnOsUzFnXUHWK2
fns1DFvOf7TRCa4kVegX+SJe0RSt7AwsZ0u/h/vjkjWgbTiJih9K1SRphBU5ravn
XY+534Qce88IPhVaZo/S9yJagZ/s27elhIwRxVKMPsIDDHfBpRkrw+ypMiVKOBDz
UmjWkeJ467DL0kQkp9dntDcQruNx0kv2a0kOPqa+kfU8pZirvBLsib/apQ2Z4037
Pb1C7wavpI2XZL43CE5fU1r8Bwl8D7P2jeL0BAcd0mhFGXfj9xY8YD+I4s/Dh4TS
w1z+HAsYiF14ltn5+PXtEwDpowb+st1ofy87R5i36xqhOpBT+57FwqMR30ZnLYBO
YFkT+yDuH/1MQWon9mdwGOhgjlsbwp4VC8B+WdKxFGtwkofIp90Aq4z3ZWes1mCM
rfzIxX1hWC/ftBubdziBho9Fq+mJgErPRWvmrPXhVVMU61rHZE6nUw0sJVw34Qxo
miJelOrmNXHN1SGuNmV/czd5NrIJekSwlcNkCR6HG1ib/QfulnFnLd47e3dMTrYt
1hPUm2iaQ6u94et/Lu5Oemb7ogiKGE1uhcwOSdgmCOoXjdMtkmr4O5gQn7Wvt//M
w+7ekgTCgX2ZSOHVvi7L4olM6zQxBGW9ucDWthTq9dex1gcYCHIa/+CTT3kJwAmb
cwUDaaAa744DUusYHpYLJkhu0vppr5pj8mr1RYpDEefUeVnSa2YT2KZB3Q9UGtDc
b+RRW1uIu17tIP0+9qmpwMa9HiMJwlxx0LwKowdsGSejBaTeBpJiSG//5ewBO3R/
AHu0Spbwwaws+cyilS4jbLoRU7ZpUGxApmKHfFlg1n7v4smJFohOqMHGHomnrvGo
b/PabfTd8QLLmOqAx1JAafGH4K6sGlL8Nc0eHtfQGPztvBAnECcaBMuJLVmnbcGi
m0mJL4wxWVeJ13rzPIN1XKK4jeNoef8mYDpnUfXQ+C9DIm0iNx3iwE8zW+5w2r9T
fOWks4cM+ZoJpAvaFMLQnH4C+Cca5OI6vitAUCaYMNE3pvn4q4iD/2YmZaBGEmph
7iHBvesmGJvGB+2oehSWpT/+KKcBY1s+rZEFiLTVH3iZENjXscR7z21OLBoBen9M
sKUMclig3q5MGF4p1YTpUgcBVu8CY+mObxh/MSJNGTt9wiL82CJwfUHVeOl6uAx1
xZj3t9U6x5ClbB19B+IzA6ekVq5wHq7tkvojko8FiaXoO+n8xWoSN6ewmT/S8Mft
2fCKkokP1GLtN0hq0YlmK0MAMFU6jAgq5hP5Uk5SsI/7JOhMghFVBu8GwpFHo5Lk
lAX3ALYyNtgC9TN3lkLtKdDYE7Ea2VVlURT9/NOtxMRptDbkzndRIIySZZqMpyTj
rFiU2/m1z6AHfmTxdpXcKjGudrnethhJ83ZpBLXCRpEQt7A7MkPIJ8rI+aGohYrL
siItDbWX9EhL+ml/yyddjcqtXbU9332VHTx9QZ/at/eSuLU1ZGVBewQafuhAYy+V
KkiryAgjrOXfNdgMqnEG6vKmhgYtfZs+9pllE0JolZwyTEXuDG7BotFwwSXOXgw+
OXCHQOTM9vySIvm4w+6WBjjNmPTvVUgl6dKRV+M6IPpJ5u+vML7N8eGOx7wL18Ok
/G82kOb270Je7L6ZhnEQY614yupA1p+7L8ixRTq5P1YsWt9WcODIWMo6KSrrBFVX
bgynYY+miTrIZhGljZPGgYPNPFjVr/zHa5brBluGIho1vjYEHqrzPaayzvHCf7kh
bWaG4Exfq5q1dPbIuVjuGQGL3Bt1uuRXRzR2zgCDTlzdksMhLwZwQ16Gj7O9mcDk
aS6ffxVjJ3zLaQB8YMAc3t87nJR1oNvjSwqq8SND7WrioIgdNDyC+Idx+rwnWSBU
vj2aeq/BWKNt2c4i4mS7/TQvnmbfLR+UttwZ5zGg+zT02Wp4k8P0mNArX+eiEFKZ
x3NbqTEWtzl7nsW/FEzWbFXciU0XpRYCVvUAwYOX5CFNUlILAPvJfoQnk9NxojPg
wZXJvDTbYGWc41OeP2E7e8BlmcycXPBOk1EboHA2HWnM7O5JaOcqoTFcsJEpftIJ
UUIBffvmDMY70spATgkTMn2cKiYFlVYxsxxsMIw8K0Zd4jcQ/ISy/yKvDHwQMsjA
RVdHdEBQiVu5LmmXW+ZYRodMwkmmYVvoZ4EopdSH+M/CXnsuiP9VCJXpa9ctXElm
zJrX5XHZUhtW1H44iKNFbII3XB8Cyoh747T0di/KukhhZsDJ4ndjDCbcf6niwoyU
TkiNztxnHgtY3IflLbT2m2EN9UgXhfsEUz4DvvWR3U/OF7OrI2tYqeq5ytF7MwHC
u9VB4OnwxaFXlzk/5ZHA4RV6AjZjVeQoLyFp/scJTp5xTmUBBRXzXD/kLJaGvHnn
2kYg7tgbYW95VzQqjIAgXzN4ORfjHtvaRxLUQRg4xAc4ogjZ8IPXUYlbxWaWzY5Z
CWv2jZAls/6Kt2UO/zqpRlRAWQs7fBwupc2HoA+5+6xepnKr2bnReiGw44vOxKyz
D8OKdeTeDNEO0wBDSLcJyyOKqsys8XWkc2e9wnAaeBzKIaK9KVwhMmoQdFFaenIA
2scYHNdJmmYT4LetWxiZcM8JvyljqEX3biF1RctPyClw/H5+L7a5zIWGwGsJ+QSi
A5+Ja51GSkW/uY+yqBD3F8lIaVW681MJ0k4hUgn0Jz6Bduz3zn8OGLMzHQHwOdMZ
vJZ37YW0r1zlaiVx94imtM2GxJ06+AsieehLSPpKSWnKSoTWMTFXWtNZH8Q8+BcE
3M//3Aluug3fyzFjWo0PitnuLdySgpccvrzv/UpmCZZqBrpCc1ez2sfqq3lzd9EK
yfwx4xdyEXxhHCq157cXb+/+zKW1ZB8Nlulx6sIvlkg1l5fi0oq8VSxLz6jZOHkH
jVykZIQb9pa6cBiAAKZXaN04I1H0VbFX5Ny+xYBfhXaHE5kRO8EZk41+kQ/LwdAs
SIbDuKoo2Fcl8nw/d5jQy8pguyzq7bxDThaDBx8UB2MANv02XNohFotWsWnA9vnx
ptLtVuh5ysL1hxt8hCnTHddICvV3FV7z3Ee64nGEw6u3kzx9wr+53BSMtzElHoAE
BXeq1mhAxoKE7ZP2jbC59kwmvyMEIZo8/OnnBugIp4QvvkBAH0/frFIRRAVOtByN
l5DTm5NaJk1ucAZNGCY0T+ZI84D/73UQmPnCCfUGSnnSEeaUR5x2VaE/WHua6bK5
MFlOf0/C5OD7zbAxuh5hzvwCVyLDG6R93mUaVrupuj8VxhMozfVnZsWIBFRAAGUa
T05QlZN+HPf6o4YLODXi3wr/Bz5bBzv/8pmWNltUbSZZtOmoAv9z6KOs6x19kQp1
vWkU+ptsFb1fDgBbRrk8B+Hcp3bf7HBDyiBKfwmToDlnD4VuN/72w7EunYJnOrK8
03W2lRbrg1ArFfCiOQfIU2BTpIIrE/DZ01TpqVnj/w+fwzBq4Jw9PaQJsFrJJiH1
WnH8MLDqF2MdbTwoUiWy3bCe7RsK24pNX/z3N82FYHFqMUpfxUnakFhmU35pUIfj
dOMHm/rSlmFm65ixchS3meK/PP6unKrSpgRylosW/q8sTseJB4LzeGrx0xJ5i42e
zAd7gpVOi2Htk/8jpybJdoM9kp6C7sfmdPFOOEDw9Wx7nj6nfMB3FMgjt1ZcdK7v
r1yTlq/17pzYhJX+9tW3cvs0EVbIy0/BP6xcHXdVKKxDNTXpHp4+HK+s1ablY+PA
5RCszRE+LK+DJoCfxQHo2gFNvoCULcmB7bdwrDUIDCa9VO5eBpXM8WuJODVo1yeD
g2CckqO3z80VExrS22T+MMIQs7huUKrckaJG2usUS7+Wl/SOLnIZZFo8SlpwBAvz
kW64uROhP/XoPEnHqFElGybpkBfaUwCAvhIWSKzSSBUN2or2YD/PEj/31epAS35D
f35WtWYkM6mQT0x3tCs4Tx+11lCUKp853zQWeyq6mO6MWVwjMsM6GapjO5Ze9dY3
8c0a8YsDS3qFeTWSau1zGrVH4+8N36vuZ2XZD6MUXnohM19cRIdHfhWCDvwhsjXh
0G7k7jEkeU3eGUIvLF3f4bX+mhiLUU7rt1hCpCUAgALpLE2b2lZXXV8CrOMHwD50
wQmp+aJHVmafjYTDExzUOHR/3TvpLE1BcBRLyTPiVvIUHmIqDbdGGdC+SfmV0OeW
RU7biHt6wZwm3ydVi+8UgLpoNeKBnzZjbAzpy9oWM9Hvpl5zSFU5Et3VCBPeZcOq
g01M/EYr4BzIe4OhApmOR6dBwkIhoiSR1UZZWpTHZYEYV8Z82aj2fXDR2myg406h
DZ5nNFuYAjFP7yC5lMSkNX3RlrU0S3rtZx/k0Qw7XQ23Fn56IIZVvkb0VYoiZkwQ
kcIn34SXbg76pGxQ7SgXkiZzVMbyxRS9isXNsrOdXX6IqwWIhujJQHOUwx5PfCss
ZyGFrn1ZyYNyxa9u5/Zw3ntS6CgjDyHDu+IOhLEVmFVC1+8hZkrSy6QoWJdjjOZG
BQwykWqUBjqLzPhgRLDatkm5W7rQoebVd4PqgTisYlPII95WKPXZCyyA4B5wAGE0
J3Xkp1zShKh8lLkbNWFuq044GvK8xYwJE808PeJbH42nGwZeNk7JPnf2wAvWr+Zr
9fmN9fFcHgfa4D3S+9Ccy7FDsYCj3dsMnxGQlj/6xk7skTHaAImt7ldNws0jNz/y
73vvGzo5FXtXYEBgnNZ95oFIAHncQpzhTh49GjzOtbiPP9toyEUhUMV++c2/+p1q
q5awE/uR2WLTSu5fZuShRw/p99CQCGrdLRgtNJjJqSSy4d4yqnkNUkT9yGysARmq
THgUxWh6SZYPHHBpzuPiqEvCslHUrvgvAy0vpwqgxj5YG98E1bOY+zybaRfkz7Wa
EowOJxRXRxiK+6M+yWGOyf6vbIRbESiZd5o7N3SsBu1oHyHfplJesX2FGvartJww
4qd/Twkmz8fJ+X8kytMuQH0mC3cxWwwOF9IUehaGuq1uX/aZrgeZ3uXGFPIRWFOD
DdgB19MILdhXKMqpKLZv22cuSzrzpY644Ty1eWG0lX9RO5zNob1sTOjWlfrqn5KQ
FJwE5k4Ea+NI55sVkWW86B0e4Wds2u4iP3v04KrYgGnNj7kXsiTFOCXbgPQSs/r5
shTDb3mqvy6SyyVHwUkUFN+zXmkyDBn/hjBh788t5ehJU4zFcokfOy+2+Mo4HDit
gy7RLMvguS9poxLKPp3YlJXeQPlEcEqySnU+0e6P6UqC4C7L0lOfFkiZnnOI6ZrY
YIdhXLrWrhIoOzE1mKxwIG62LkKIxfKDbsANQyASbeFuu9K1DHar9zu3uUg+YLl2
8iBHfs5ycxyYJkKN2rAhrbPLnsQ6BxymzdDwuXIaqMDYoK6RxSb34NCX4l3X4bWY
F0Qybcf2YDMC7adzT8QTZ2GhtJMcacQgwBJtuI0F7/O36b5LYNCT2ww4075M8m8l
sGi/2PQYgsW9oGPWLpuqHlpGrTfzgGQSoas545iS4Eye/afCZTQWlQdY7ixVo+wE
nEtt3nVixGzbYPCyg1771PriawhhPEdLR0Wwfs3CLRzzNzKpLWzMhjYykTaDEMQY
q/NYWH3tvG4MsMpZdFZrMyfwKs45qNjWZBeu0tFOnqaNLjyKX4+D/vPSuWKZ+MOy
rzj8GnoeusZWugt9Vo6TCz0f4TRe2HWH8jDCd+zZqbjLNgD1KnYR7WPZ1ZbOxrrZ
Z5yctBRtc0UP+s+3PHr4CBftCIo7HaTFRAMgQV2k4KwqzB+5V6Gt8LaKVV7Nrnjm
Z6xr0b4hutffEp8Ftc0fe9y3j4VTcbwGa/WpT+uGE8N7w6UGr4DP5WGjvV6hikL7
i3vN5PYWBImpu3V3ty1SaDBRLpqIJl6PzyXqfexr0qox14rlGgDm3jGFxO3tpL1S
FqkiPm/UxJ0wxD/pKBJcE1f6c31wEj8xqSb8zjbIeLB3pNGGmT2M7bxjIT/tDdZ2
PTItOF9il2/EBXn9QszEvlHqR/oNz8hd54ajqxrcWsl9w45NO5WJ/Xa8z2m9RtAV
oJ3HmR2xB9w7nvtILLa93NZOoJoVHllGgkhVgjQnzycZtp6ArBs8LGuKHUxXXpqR
nCVvjdJLbHiX2JujzZpaPt4zxujjIYLBQnNA0wdUqAV8rfACzv9Zi+J1vZ5KouAU
3QxXQtH4LmNaGvJXy5nhCL4GKI10jUFXUh7ovuiuTJyzD4bP8oxO3Nkcrizo6Kbr
SuVQYqXIjAeKTeiiRxiSNv07wO4T0HCF4wyMt1hzgAXo+XIzYUgM9SLdpHSzvsSa
a1kIPxSrbRQFlSgjfCwD7fbs7Rd0HgiPpzokysvFIIw442kn1wuGQfszDlBuZ8/n
wL8QK4Nu5+/XHExWDYoRWrsuNMRmkgX2k7mrGtVVphH0QM2tSUd6LG36lf43QSZo
ViAUiWdSa1XOzKuOOVjocOcLGmL8phXzv+P2IcR/5wdJfwGZjvKIoUHYBBkPUI2Q
MgbnBWkK4qhdP3Zl/laoDhGOecQ5T04u4n756qkIFfz6FB0ScwW5ZCezd9BotEpj
kX/NfC6n1ZDFrqBeMrX40FTIaSdVFLhWvD9BobuS31AAJFtMuoSK7wtqk0fUDPlw
1yCgsnshIG+YyI2Ftk936CcjENaOBHQ2IwN5C0GJmwlcZv2A8lRBlbVV/N5b5b8b
JIQqF3a1MgEBTJ/WJL3Rmj6YOECE5ymjXJnkjzpFDOtF2XJfMv5g1ejO6i6XGSVR
SHFo4Kh9quVP6K7wIpxHEYnCoAfzi6II+7XsgEoe20+F2G3kOMjsjqOOQCwzFLJs
EfluWYvSxsi3Egyt4KVZceQuapF3K/oSrc/w/7BTq/J8+XCGVZJBV1xNQnTxnmnM
ry207o15iLWoCYKpeTsIGnytFIBOMl+5JkCU4ATkjRLrCRZE4sjzfOG9OJWWsd33
fLL00N2gG/rRMEnxzvkfZnym4c5jP+3lJ/0nCWaHOIeaIELHlY74D4buf3Psgzx6
/67YqkLTG5opZfpbpM46kr6RgODB/6Qor/nWK9nVTLloIqgQXpDsl5De4+wNOOqf
s03tDmjy2Nxd2nAWkVbV8o/FtOyQFwKSVVIAcP3fEYq8anSH0FoJG5K86QE0lmRi
/mf9aV+XpkS1QVuc2k0Q3l00NhNpzlNkjc5v9Pw9ZvQ0YvlMMxGCUUKtxodXYfIQ
yedc5zzglV/C6/LdKYtPQEwdqv3QDBObixmRKJc8J5HgYsJJNv5wYqxGZaLz146C
RieIAzSm/ccgElWOgDk73uiNsBOdIYS2YX7/xbXy8lci4ivjcLZtWhh3EPodHad+
2+pu1HdvcObp9NB/KlhKGCidm8uQ/6PBhFcgKZsIC30k0prO8x+03CkIFt6YheSm
apZczkWEpSH+L5HMDBgt6VSodwqZwYria5M9FXxsGorRJgq0yYYlRFRxVTb+97Ah
bt+nviAYpI7AQhd1zDUKKmkIEinDLUoKP9btq7dRHO6OcgtT5sGIR/HU66gH6hMo
pCmTpTF2tdrdev4/7J8odvJvMMEl37ACou1nRO22iqTWPI/swI8bn3HZklZIf5Hm
2qcJ+FQaeDdE3E9WUcW5IUmuydB/EmUtow538al9Kb2FhTuLPQFeRHNPFmdUnN49
GV+XRISpB/h6HZXlgCJjxvHAwSRHgU+dEfS6DfOzm9r6Nxj7yTbJKObr/rRx4Mij
88yegPIrtJ8C8f8ca1EvYnMQiBiQz0kW5YHtKKrgeNErV2hzMu7ihdnidomfGCAH
yfauoUsy5RVhkwXtBCwkCWXEP3uGvL/LY7y9jGaUrMx9Kfu9nTyeaPUP3ra+juN/
0jJbXO4Ly6r6+cm3H2jEdGLd2OlBVWzrC4gAZJlbSe461NNCnknh8okaXDsDas0D
T8w7rxiP6cQLDywHrVtN43p8sF35VflC0MoGcQp359CU2VoC819gzaLcDM24z3CE
8y6yFaskSMX+wfSab6p3ghrcwgcZ9FUpW+fItuxUQvrnTypBZN0OPyLvl9oq+ECT
AP+bxoq9ZBdKuJTPg9u8VFMrE3LY7ZPVmJE+PJOGvdJZXu4yPrCU3v1jmb6xD/+7
ORLpSr7hoPA2vy7qjr/KmbNc2+iAA8kgZuDIGHxuAHagADKpfuUcsc+mtoNn245F
kAs8iYdlMyIR27bjZIX/PqgscnoVE5xY2j0dvZ3ZDQ8ZRLptKjjrNRJ/4Ss5gEmM
J17iICjBJI9xNr9o3EpQl2aRdStXyipfIvXRI6Kbz7VaqqHUlpGrssLMXuDRcURe
SjM/wcAyxwdaV92lW7ZRWDix1jSyfJwswAC97QWVGVorX8pCr823iMdg+VGM9+wt
RSf0KhOMvpfu5DsdMjabMp1JakW8oOApQ6UbS/oNw84EE/tI3TP2WzNYSCu2QfJ/
NDGQw+UgTCNFyrdbu76+OHhkQyOpV0QEucLaqyEm/XCF+6Kamc1Rg5bn0jXoMXh9
dIfgY8t7gsZGNnJ6F57FHmkQjcMUmdi8XMS+R+/dlpHM2CCnXGHR1ODDrACHkREZ
bhxm4JMQ/tspV6AzvQmRG+F2p+YHdOxhkq9BHwWqtRxYNEefcsseM4FQnanWWoXe
N4p0tyz8M6TmQq7B0LAgIthu6eHdBka8C/NhgbDa9Xr1RKCsTOsEpIfbLoq0r53s
0Qc/sPj2gpxYvnm15C5SXrtrY3y03WMtm4aQ5gpicuZMICTBaMaIYlaGzzEyAjEr
AzixzFZWRxEFfFPVGqR4phFaqKyZFAAobjYXBsuRaLQblaKwmxA0h3Bf00cPNDVW
b4RU4ZyTlFu75iPdPFAHKQDrugkqveGlyWB7e2VvyywEyYlJFg5pP/KAA5Gxk8ID
ZxjGGQzrDEonxPWjqa72GsnmNfk67n9H9/5oEMnQUfsUUzEVThwq+guJNZp2Rk1G
XbTv8XiqCaZCns02Fv9n6Uh8ooYTQRKEgXaEtoR4KYtchxtueS9xCSLeM37bCWyJ
xVX1j3CxfN6xCZ7cJKko9bvJ3ZhhCBdU0sI/1P2i6Au3qcyUOfrpLc0FM1+r2L/4
X8yuwO+ABpYni39t5kU1BHwa+wws3fxcoOXMSSv68mOdyo5fPL66d2uU7g/uXqbU
gDJaF2s7M20jiUfr2CEqHgNsjh2fnEbF+jcSHMQ3A4z0NF4Kmo9yACJLhi7vj3Rc
2rLepiIdYNTK/Vc620ERWLk9jrApRRrFBDdDkUsFlxBKYJI4SO4mLOYfpeqZkehI
yD0OJzV2dUfWRMqZuA0eca+3PY/NtL4aM06w4qpwYFEwVv2YUP7LO6KY8/fSf6Cg
Z96EtY1qemQ4+6yAx4hCFP3EkdDkbyRUI/XFSsTPcScNSSkC3Cbh3YmXWTfwB9Z4
BhSWaeVE4sZKebL80+l/I2+5JsfFUF93a5oDXzY7DY2ASkofiPWsvAzjcItA4HZE
jA4dcC5chL3GEWaTUx7fezmnlPDT8M5oLnQr5stVWLgEe/ME8gYjqB63dPSO81Uq
Vu+vBbVjAQHbQF3r8OVi2JO5vgWuniXmAU4YeoX2ASkFaieCaVzNdsTw/29k5ogJ
/6CNg5rMsrh0H+h6Qw4Sc53Dgmgi4Ez/SeTHpYo9/YrN9ca3kY1kOKuzS2UxPLSi
q8SzFcTaXwXk4ucTxpshCeY8pJ1LuaVOxxfM1qukYUdsVQwgmb+uk+O4ehSVoqTh
2kp2bJbreSAp56r/XE5VF5W62h/F4WwwMLgAHQOnAMR4NB2YSLRLsDHk+4EZKiLG
6jHMd7Skpb9ixJhqRptS75TCfsy3cwNHRqcpigkm2ZCBWdtj2v7v63X4TVvJIYqf
jAT8pYgE7aKCxDQu641/K6Md4f3Y7WxYA6nF53cDOsgQi7FIFGu4B9pGky4Kqn6V
R8qQPIyNEfV0sMEaxYQiAk57YzJk9hewjWxUI27o3mh32JnTlj8c9KfTVPz5Bs34
mSZtXGDnKXhXpUjheGm15NyVIXAFUCZZERIvgYaPfwpz0UU9CtEWjnjTUbNV0TQU
uGPEtomM4lnYwEK6t9yCmRNKlyV9bTQ11j0vcXTrh+OPuX4u+fN6uv/dH0RDV3Eg
MtWt25jBgA5Wkfko/ej3fg0OXKiZXGezm5nS6+FkeNmBVRUZqNP3Ud1JjWkGbg4J
C9K60rR9GHOBOWCiUh4igIUOs/lYzgNWtsaG+ZXdojN3ax1JU51sy9q/GceO9GT+
eAFwR3FbChZxPgE/KHqw5bPGdMMh4GvnGJRRKjo8NxmW29qaDNwNQshh/Cp4L6jf
gZ3G1756A7PjxD/TFM4gBu/Y5vABuYyglk7vgDweXolijpHm69vMbldDrmwa+YHX
zeNaWEX3AggqgqSS/kVUhOiCH8c6psHwJufgzfdPDTesu/Jx7Zx6Z7+AnTAYwXBw
ihKCbWEh+cbAOVV2d63Jw0xSXQmmc3H5SkbKucy5wb+383QyWTNpph9WlsYInuTi
5T1Ardle4XiCXwypk41jUhqUXBcVWMV8HHejSoZGYUYu9HYxcbcIIXXXCnh3skcq
Z4aCuNVfAMUAWzPz8VWTIFIi3K4GzoX/l0Z7g3lDLJ6wmhjap9vE1AL53/gVpM++
FI8HOzPSKjWzgm1HHBSuvQtOOpQv4nZuq1HW0Vs7EhAAnYMwiH5O+NZoggi2QkY8
DHknskinsMjoOjja/M5CYNUgPJMyGNynjrat+LZsp494rH5uOWpXre19lE8pmLOn
IbtdlyoGp7F9CplJcACLWep/QOtMAyV2VnvP+KaoUZi68IjtTU2+iHjdTDCiYUIp
O+XDXOPd6RLBxo1Av0KiJVkl9dHcYOsJ/xu5qrtR+yvBlelAoiEOkZRnhokfY0vZ
LiwQP+lr2BO94VhUNzVOvxsJias5biLg1dBXzqgUI+r+aEhSve4YBml7r1yUyApZ
3SdJdXBaVtAae82czDOW+3IpnQ1+fwLWL+7kAtphQBfjMbt1garkK5WgL0jL+3Dc
JEqwzwqHq9IIhc0HAlG0cb4Z2u2TAfb6A7cumDDhp/zHrYwL31Y8zkrFcKBDUubX
bkXJe9aDqYutMIXB3128j6P/5Jgsj46RYu2L7/b8lT8VD3xRIug9e9KbNwsnk3bD
PT/JIYA6XSRM6qQRtMvHnQ==
`pragma protect end_protected
