// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:46 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Xb4+pTJhP2ZCIaiSFspf9/e5YY3IZI756ck/Nk/+AYg4RK/0VvxymdUgpnQdywVt
7mUV5yihIxklb00yrQ+GG+/mXzoyjK+Tny9qnvQS43BMqLcpPrBctqleC5FdsV2P
VzGKat1ORjxo7LDn7kbv56m/WwJ/M2X/kkBSwHjchdk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 32448)
yfN7DGRF5b5nbDy9LEo8FgmAy6vLO6X2kcvC8736u2qrHjevjXr7VbYz1hUMd44j
Ko0kZd8nW6YQ0L51k4NL9fb7u+n+1V6xmNUXCbZ9pe06ng6ceLL1piNvhr4q+Zez
yU6dpJR7Xx8J8g+7oh4OKgyfx33FKtTDjKSd9uDoeFHdnpFvdn+5XY0oLPJHl1Q/
6UMRpZwkf275aKESNL1GsC8I2sGQ7GyNns2Z9W++JmrvMht4ZSfkuv3P38/QZOeC
OgxkI5Q8OhmBCmCoGWi+lzXsndmLdrta2L4ZGOeZ9n2i0Ie3XGKFxtCpPaGUdCfx
Bx4qkCuaqg+RhnTutvfABJIxicwWeUZNKoCKjpXnnQL37XOHX7PPJ4TeNVi+6/O6
lOfSjEaYJDiIoMvHmVGhLzdspyzaRrowOdxlqVHH+HFOYGwp1XcSpOP17Q3EoV7V
g91bILR6/jPaCnQLvj/m75mguRmRolejKFAIiCNlRcyg3QLe8+PvOh1DX4FWdLQh
O1/cnQ1Ku7XETEIO3mdRE3ejWVxROXrFsLnzd5YNUzVgShuM6YohmvdHlyz1c2Om
zvQrpZ2F6LZm0m4a57IyfIJWKdKmUkASZTli+jXIQYG9f/oQwo17jr29WLHORYhe
bQ0e/c2u8GuDGzgGX/6GCnd0WZtCaXHizWAj/WUJXJyUP2wCRbMYEiekZhMPTM36
ex3sIIC1IwUb+OE6Pofdt72a3kBvIyPeQ3FsXuMfYhZcnXxM76ZlQabrCNbiiqDP
zDpxQbFNZcLGeKgpFi0bLhH6o7FTtServBr/X0M0qrrWMBxDKHDZAD3ejelmmAdB
DFce/Wg9SNH4RggaldYqySsC5PFPo9KIZGJ2WfdHNA1VXb0RBRZhIVEbDnM94M0y
fHBOMdLYUV/nzhSuFVIO+KvyWZxWr30s+nJUAl+SBPZF/dWpDNIME59WfZBiwM1r
IdL3YejD7hPebwXccg68msHqsP+UU0V+e2I3gjy8lWIshlfTusk00KOLBPYWQ9Fc
yaYAtgjzoBQEEopSxezRekO/I3jAtBUGM359xKNZ4i78SX3vHzYO/D2l4RZTvs1H
6ztplH3HvTzvFIR8i+gHyKedfghK9FU/UcsxQV2MK4FENlxE5iHcONkKGYpwnZvt
gntzweRWhGNHoRgljEYSSwboH3hobF8US2wv083rCN/orPiCs/19ZSi3tV4B2O+X
s3xZVy1Raqa7Nh3DDFfPqCCT5Tl2fy+d0zvFemrLc6D9rUPDry6hWy1WxtUIH9Qd
nZPWySVJfVUau8Hhejc9XM2TJw3lgyBoG4I+zkLsuWCmTcUKeu17vMWdC0r5d+Uj
5ARdqlCnPBNrIgI7K68sXnISD7Zb3N8J+mvs+4KHUXATDt3zrezRou90ZXN7REyb
CLrTniJqjRyFSTirb8AzHd+PuXm+NCTY+fiyJiF9cG1qf9zCo/HSRnBCkxkqrFFK
Vcn5JiegYdnhXFobXVxiFl0H/P8kynoIgBNFAhKPXRABmIL8YGBmz3moPKqD8dX/
ge6cEcca3EXrlnT9WUomRskxSc5kfOM7VOPYaJXW6BSBThEoYYV2qShGHInBUC65
8k/KtBmMV1vWEwB+3NXWSY51Xc2Y/XFTPOGAkuT9Hpul8vq0JlRViqXqhdfCUECO
HTrm55LfMsMvEdcUvGNZeqqY1CIEb8HaC7Ut3mC2vzsRMTXdlVv5Tw7YXO7b6WlP
MMKh/4NiAG942/5EN3/zkw47pD8Qy2IZhBDKgacmX7tDU4JWbGYRX54XI9lWPEvq
PJZ5buaMbJz+1twc7eZm6dZSolOHFoeypQ6+BaWbgvlLYMPs2kzEVOxHxI3NGIRb
QDfiGIN8HsNcs5sp1aQTYZqyAkdWc8OXrTdAooI5x9WUbj7trRp2gA4vA68dhQZd
aHQLX7w/4X24smbSB0IBYrbhiOWCnTgD6yLPKit0KHa8wiYaJz+itre6p4HxAzXH
00wEUlePbw17pJbnLxhI35C7/Wqf3k181101saiSID1RnJ3VxHwmwRpffZthj+Jf
ZCBmdLWp6fRkLzZdQkkeq/UundZA78o9V0lM7CIFFIaYUicmwiCePRxJVK7G3dW4
eujbly/0x0JdZ+syfmHISu764TKbg23jh/RsE3LIg4n9LJH7faNqOy9jsSiIIlNX
dD1nE8FFLJ5iEUMdtEGc/wEI+eyghhtXXD6PN+ee0SDuUuejJ9kCN001/rkYC0Mk
stflVfYIN+E4vGeBX8PnyE8z/NMNTjvd3bCBa94FpbajnMXflK2Nm8ea7MMqkh3Z
IVC89rI4yvISJ1st8Q+zrsKArtLjoltlUsXNld/aHPH0rSdhRsYfxb6ImzE32GSO
VjeIRW1OdHzeOiHBaQTS+ZwNbipP6Sub5acXFp8/55Iy66DtzZQ3DT6d+j16pLcS
J1QnSN70o2LpU/2Ca6iCW67vo92hKyN6LJNnMHHXM/UICAPPaYZ9PJ/cH4/hQwfc
WtYRRoPR167DCWKnOQ+ZQMzzCo0vk2/+ZKCkQ6GtnRCuaX4kPqo9t0Ljo7KMa48d
hN0/9AdNJ+z7YlAPcTtCKO+FLShO5r7PnSNwx/6eH8F8ENNh0SphU+IBs8SYL00d
UdjZAMHuiJJVHea7bOkrALUF2zPmj9s9ycnlSv5x2kyLP0EzNOeY66f0Qbejz9Tu
jm5IK8pNUR5eJlxGOGUCETdMVQ/jenCS/MDrrfzcNF43EUJYCxVR8s5CrgPfTxWI
bMiZdTyEDVyXk8OH7715wzP5QJoRGiY9JNuwtNSInBnNqwugVKXIsSBs8+C/Vl/g
Fb1F9f5rUBPmfm1/G6yv6zHYpTmoIIEPJUWsX2brqFD44b/83hPKhvKSLMQaE2P2
I90SKouEuSAJr5370MXwbRc2URsvvPkwbWxSjo0cJ65eFYyuEKe2aKXrGmHUG4Ug
cYsd1VIsVPVcE0Pb+OGwbtsFIi1++J3I7/l0LeqTbLjr0ReoiHEv40fMjfCZmLOE
RYGgjuu+N+6vkBKeCJyYotBciGj1pRIxgWIQeU0L6QCFxqrrglOZnz+Sj9Ms3zqw
XAd84svZZWuHRU3R0MCfd3+BB5tlt3EbECu6NDchHcbZeeFHh6uCZjWElz8DfpWy
7oy67jL1rPxlVszRWBFJyR4QN7Fr9JUNjdPjT5A/x4RQzMydY4sM9yRI8r94JRam
w16mr8QmV6eQNylg/LRz5HthPwseiAQml5rroKCdiTzsRN+lZOQYoh4ZOvg06yKX
N3GWNU481WgoNRC8+I8Owr0PPd4xGFNEaQnk1Pi8b+VWmzimVwt2bF7OWxsJV2R7
2q7doBPyGNSZlvYxlNU6ILn43is649IHxxtxyXB+cXrtnTcdwYKX2q8coAWB99mY
NRKp0TySH4CD/EI6qaAa2hIlw+UEtXdLqD0m5w/sRZaOfpdd0T4Jc4oaCgX2yruk
7fTLKAGzscsCo+BwslbF5Ve/ltoRZBG9VDamJPA6TVE+B9R9Q7E4WCrOHSjTFv5d
WlJ6bzT/DE9kZC9bzuxMxJC+bvD9umgihTguqTk+ptZNI+iaNjlWu7qE5908P86j
lS90WMiAOMOYtgijp7GoWghx/Zl+3EbIEASCGpx110PslDeJIR9KkyIK1NQSK5fX
9hXjblMSXtJDclEkuqLmDReX3msot+VMxHe7aFY4Swvj3YcwFMc8EsuiNvifxnqH
aiV9NjKgYdzIwt+8nzGFeggJba08JlMjp/K1vVH0HhSa9V/0Pf1GHf4My8OGjoR8
u/THctXRj6nPuWCGzY0h6TDfn1OZ66iVMpYs17UwL7j+3n3OV9aaQmNt4CRfWyVC
xOTT40Grj8xu2lhFuNLIBQscU7Nn9aygpXVZLIc8/DF8kvby1eL58UIoRe6OOBTa
ERihqL9EdRKdO57kjbN6XH6x7lVNUHjbdaoIMy2YjRvRs9l8PfZ6FSqy3gkiPuhw
+gln5idiZoAZbY+Gp898CcQ8Liae8GWNUtLDMMS7mOFokxQAJYgj7Z42a3RIKbyO
dbl5SfhMxP3ROfOZ1cA6Q1p65qPQ4cBk/f7ACTyzyJX0cGbFH+kbLwVWKXspjSan
Ca8GUpu/lWtGAvJ2k8RPcb77SjJ07QPt62Yep5kCl/iCljiy4frxydjJ+1m/p7N5
7OHM9gN+HQTeSsB8nwDMlYYfjVv/stXGBe9KR5+QLpi5ahatVRvcTuvlmFgd4c9S
XNTbkx5AjI77QbAEqtUcWfUR43WOdc3Y3xRbUe8fRineV7qAynNXiaX7mgBtNReI
lAxAf09+p9q9SJYxUhnyQajT+4drptVIrHccoEpRFV9aJq3ymEiwpsOK5eI/UMnP
uFotoX3tzqAz6lzrFsl24cWoqPY9mZ+XBd9YA5y+wXvtGyyga1LUgSThTU9yovHT
8cwShyTZDqP2z9ruup3XEE4gNNpqumDRhgY+puzW4lUjcypNbDyd1usnYVFK4yi1
ZfmYsAJqR0EZ8cOumIBfPmLyPOTQYIu+ca3cZIhHfghgixZPreBQfYJGEbSmoH0b
5Yeu59vz8bUlUtGRmu0GKNgW2T0EZPXyDiCL+LNpQn0YxozDPHbMa6UI6zqSEAgS
m0bp2lce+tR6qttqsLiKkWcWvmmHG/anjvW0/OsA1Nt7MxyoSNyeT/sgN58INHuI
9EGr/Tes4tO99tKb6mxMDT1K1dnJ0COOq6WgzwYQsCqf5jUHtAcPxwVngrdm2p6y
PraNm/lRUAYxC1FLIyhen1kp5lNPBjA5npeFCv4CPrlRjTRdhmJobDLYM1Bj99P6
y+lWFpFmgI/JeGO9sFZcMNs1HEgL3oyjDhkVRnytvKzWxwIQcL0vLdhfZPZKMpqZ
Lodhzj2iQwG8HAqzg5ZPGeyiQJHQ2A9IYyLWiW8zutD4yG/ANEakbyRonkKFS1Gg
PGnyqK3UqR/Yru7vF3JYLuIKC8PuHAOHHcGVUOn7e4ZW+syoLfm5JXcxNl7jDI/t
GswNmudeIDKLsmHYOQASiDbcuBjmFOS5kqf5gk8gT1QRg2B2xxmAEQrQh3UeIPVd
zmIYfo8Y+V24D1qHliGoesp4AvfwOc1j7UpcD2zLn7gDDwMa4LfLksfRj1B1/Xps
li5MJHpD2Pis5E42n6H4JUiPTCRncjyLpLC4gvGb8U7vDdYgay7YlT+YdEo8oFcq
bTsmS1835/LOrLS8c2D+6Db4/qi8cMzKKmlmfmUSuCZgzDUxeC1hOxMbdjrf27J2
EmWs4HtlP1bJfcEIPMbhin88Bk0hdevxJoq+Vj4cSkw7DVOxKD3Ova0N+pf1yIbg
DG/hePf0IICCiaqCxFJ3U92PrTAafrorUGPt9NYMjimSLPxvhVtUgrBGCoUiK8sP
V5L0n2+Stn76veqS7g8GRaxz6Cw2dmoV8Vagn7XVkRPk02TJTa+FIB89nz9QKE0C
LhOuVg5jIQG77/e6zdp7Kp8aFsMVnsoIYcTFNjMeKKI/LIT37OZ3gZV3wJBCSpOw
IBtxhiPJ3ZkWByfZDZDqg4EhUlGTADPxg1KNcz1ZIDVGtUMjMh0ji9DxVyhFeKsK
J1MLDua1Jv+rszx8/oanibIWoeF/Bq2vPuHobqyp7kFTh1DL+9uu2xRHCsELfdAE
aaV0L8HcnCUwQMTQVMC47rY8ZkmOd5IXnn+exEbqHCgdqk6oSEeBbeb78ZpQk4tW
sytl5O2fbw3ZrVleoYeLmnd54ipeXCz5dp+XIJVh+flTfywOBr3YaapUT8X9y1G9
LcK9V6V72EtESZE5u8kdC9j/XLG3Ubkdxrd+sdSoB/GdLTgFA2RERVbf+hTxazse
mIqezJ2woc2O/NmGQiU1/8LWrJSxNM1NNU1nk9Bj2nPhI08yGpDGkEYu8Qoynx0u
VXRt3GzcqNJAbfEh4cr2azteH40LSC9MsoLdc1f9m5InNHFD+qhvv/oTTbDUdv25
CwWp6r6T8GuqXS05iLw7Vp1PqM1nHWphop4QJaLuln60kC2EQqdImctmVtbKk5o/
PtVtH2uXMZK1T6yL0cVeunnxTh3LV53MV7atF0A1/e6DxM1wXTZK26z7WbzN7adU
rjv4nulAM8GXgbSakEde4B5/2pgO6Tb4KbPv9tYpgelb4HAqDGVt4NPLbIW967Yu
5zTbF1SRmgu1Os8Bbatgb5EFa7xHqH9arZYgjFXDdLCe2xLDIUFb/ivC5Usb3zGK
D438yAwxhkqFGYj8veMNN5XxMsqshM9prQNGrEmHPQkvkjEqCgH8n3lvcAaJGlYA
TzURUFpwsE4hTdTh0fIBzieRJ8Ne4ivXhBGP7P4OBKndF/VKhmxpReTVToAsXy1L
WXMsBU4bJ0YYMwIIj1UKhQgE6YpMWZ8B68TPNhDTl1hN9724uG1c6mA37SY0Bo7A
U/8jj7O8HMIKSBJK06xe/0MNuf1ocebEREr1EEWA/N+afuMJVfc8whKqMRxIHSdQ
S002KYCFnvWkEFfNuMo+DUcN9s1Pu0NaehnCYM9kVt9VIRdSUMh5Bm1U78cCfb3y
Tj3pZWWsqICzIak6MvQ51W/hmZbmbzRgkKRPzDQMe+9kcL4f8VKe2wDmVXaMxnsE
eNBN9ZidtoX110bQNzDaiK85e3aoevze3RRC/U8PEsBwHpCmtpMxgMeHk4kpS0ql
cY0U+FiOA8RZ8vycInYaKrZO2y2IqnN/27Muhr2psojXCAG1OjF+WIpteyJZ3gdE
aaFa4mh+7L9JH9JARx+CyMWPFX3iCnDG+rDzpa/E4pycDBsN4Ydt8TxlANy5AJHc
aNa5OXTKkrxg1dEyD+zlcAYXQ/ppOol6nURmEwXwykPA0Xc26yQODzE+dXuv/XbI
GUNs9kHfMh+8DIh2Tmk4aYmJRvtY0hhaYo7drkcOYJsttdhRyd5hy5x1Ai2kfsXG
HP5e1Mc/dPiIPAcbV1PiVzuCkQTkTzPzZKh6cNAB8sZ6mLszE4wjami5Y9MzAPu8
GFEciZR1Us1f4vLpEavXc4mGCUZ6ZsKaS9+8NzGFyfaK8b2lq8983EyNjBsYTDtN
a8sT8EohX8QPYyEJQ69zV+CIRHUvI4sBCOkLvEefwlZHr4hoN/oHu/AZrGZpTzFm
5tz8PW9qCiPattnjGEMG0Zfm2Y5fRFyJeOKhlknU5jDM8eHeQ7etE7NAlIgag6L9
2ZKZMr9VtUqU/OL5GzrRCHUkdmeUzQgAf6n2ivc/Q57yEnP/otI/c6Q1FztvKinB
hMT9cUXofXPuUYMhag0EMXqnpNee7VH0eSQ0RHR3AxCKeYoJXh7qoL6DbK4ycHHO
gEYisFDlkMM+yexd2HlA2Fau2SyEVZQZP4PClKgI2xvkhTbwzy4iHG969ok4bG38
cxQHSss3IiBXmJAXEu9scQmJuYNiQQnFkrzKmBJK05eihXTLtJ+eAOOdN6n2oj1j
hGEcMO/yEj1KWXpVL88ahhOdMlrQPRPWNGoj6iJl0tGC6jpnPUnHhAseW3D/fvcg
BdORrhKSw48J/tmtdIiEjmpSYub4P7Zb4aElaVRbHcAmNbZYizJvDFUYxvoraf3+
QpB9W0KKcPPHrdEY5k1qmyT4fiLgqmb+lmSPRexzPp6ZomOQYE22o/cCpRTCJ6Ic
vJVqikH2nXwPkZBdf21NOTZC/xinyJfD/D8sg2mP9TxTuHrEU75gAXXtmihG44SO
JUSSDJy26HTID24LS2wiKwXs2KVagWT9iHUHbJT3UR6Pq335hfnMJq6MqCP7XhUS
ZpVmMJj78XHF4bFrr70lYpqx0NxXoqVHj6yxf3iUZQKRNxiYRiuCNO0rYFPcnsY3
oxasln5gBJfn0pNZReF4KrU1I7kaB13mMUjFDJQpx/eEfdPCoUDKdCyBm6IRIbJS
b2a/2MrOeqQ/hNtX+XyeRnH35unigPhZnPnL4uCQDreS42jao8d0ekCjHihSKlJf
odgea2USuMzh4r3JQjBKYCo7vL9CfEqrH2ZVoEoEbt0ZAxR4CD9TKP2118t7Uh37
7XK+nGFg/xU10dovp2c3EegNrGaSz+zh31Tr62bVG1NdP3lDvMmFGcqHYUJMAjJ2
tJiBIir5AmusQFNrC0fkulgP/DdcJlJ1h65cXm7qUtNpcd1TzfniDvZGnkHsZH8F
+/merfsk2yrs8E1svkd4tf2DzXAYsF+Qp4wjfdPpaEjQyGFcY+J6aOXUHNN5nGUq
q/txCVqrk5vTBeyPWzPuB7S3DSMxmqcOqwz7tJ3JxRv1oAt7ikTRIaZ1GsTiaioY
wegWoUgYP3TgnvPZWbJCXykHwvVph6075W/Lm1oqiD5aii+lrjGeJ6OrPVAZIQ62
FN0Lke/Z9dGXEOvTLy5jl8RnbwUeFOuPwZk2ZG23zFPU5+PreTwPnbC0/36mFLi4
UP6ePlkxOSlUEDwZ7RYlzzA8Ev+LCtWPLsrgsWYtM0bL8QOKlHleQgZgwrDdKmY3
yBj5dhGo5VDH9W2kiC1Xdhu8Vqx5/0VoP30/WQ68LlJYxsvFhwPS69nWoeMnlf7C
bU++V0wT5kKAEEzoFKuydnWR6VnKGL3OlkZiVegtxI9iCJT0s901emnWQOn0ghDG
tPCRrGfnDa2ONPACCd+kkI/+qC1mdJSzJJrcS9ZmjOI0r2sdvd0Vz+aUoTawo+ej
3tcxvOtswksZm/KV9whh4I9wREhhjAi+a1Ay2u6ZiaTuigCm/IiDPP/MxuoMKNuV
t3P/6XZnu1w+FcUwJ+eGoFXDuus8gjLpOseLLFqSmBL8YDw2qwHJlUXqMnDlxlF7
VPupJ8rhJiWJOKecu9DnJMBBi9HfxKkKyBk2unYxpGOSKx5BAwz/RX0YV93jRKC/
RfTo39GFdgg2Lzh6ojSfgh+OeekgVsp807TyWytKE3GTILI+/F40W0nCaw4AsqhH
VNwzKW6Y7cITuTBQXiE0LIvKpwC0TOEu3bWiBfVY4hXndzqFdkXix4uWAaJV8rN8
T0JdjPAh9XqxVpZi/OXQehEqanSA03nSihDhXe1H8f/P7w/UoD37aRNgFNXaswtP
1GPFdNecOXJw1LhStKvSOwr++4OlxdBbts6XwBMAf/fiSgVfd24tRBOCrkZ+eSrp
RAsGeUrs3Qb8/3bNzvruO52374PThqUTjlr2ihOwUQamfvh44tFgpT0k2fvUDJK+
f7UBiCNCYltV7eup3jmCE7vrN7fBxS9BcGSMJl719tzDlEpN/ZSVAmyEyhffR4mO
FoMqrcQNOUT+ee4cDSnYBUcYP9IO0qYBySlE/9u+dThbhMVibWxuWUQYXezj8YJW
3978gpYrgjv4d/ekF7hwkSPUB9Prizh8kcXl9CIWdgLL7YkHvXPnhd0t7Xx4mT8T
EH/1K2md9qBuShTMnJclHs+5Iy/J8fGzM+YsJFJBv8L9gaYSozVwN/X5xtacfoji
IB6o0J1s6JUNSA+IlqMSxVkM1e3Mak1bZfxnodFhxxy0DVty6mWrtqL9ph8LLuW+
0reGkgF9LFCV1IZa+/dh921z3I4ao4Jro4Or1LJWD9mKszp6+uEWvrjtkN+v0rAr
bMyEwuMqaY/zJQk1Z39leAxuXovCMeRWN5y0TjLV6Oowq56jTiSv52RM0dwPu09z
ghLQ8nxzTBoTzAwua4F/BPYEO+a52fGg5oW6ggW2Yr5TFAIiRgud+fGXScmInqto
6ay+ORjp1W/ujpttBV676e2O2HKwqtbBBGfvuUlz0Y6yY4I554zjYDW/jp3OVfnh
ZtSCxIZb2usznGjMmYUhTWOH6ii8EcZsnbqpT2nk6gbd3A+bN3v2ARsJy65p4qok
onL8rzJMJRRU1t+ZC0Smv9aeahs83fDjNN6BIApXuSFEzLBqzOZs0H2WL2qCG9Hw
m3QgWBpyb98PkgqRhZNetckoPy9RzEJJmGS14RSE1RbSyaMCNpz7W/YibylZduCF
4bWLl08dZk3UCjtUuITSvjrDozQu69MHO+MiDDB2yyNRLvIQrJIeXfgOzJ5DXUPM
olLDKCQYrervvunRW7L4SZykhqMRc4q75mrtHWSvKOkhY6RgY8xuJwKF9C8mSuay
ovl86Q76zARQlChxj/SYX5XlaBr+QflMPjnxHtdkrjUr/ML2+zJAhtIoZ/VeIaUX
K4fp8fDbcehNDIi8EetaBQ9W4ouFqXgRurjjqpLndkuoyx/yEeW0JVYXMM0V+Gpd
UB1w6hrumoR9V9tpeJlJdfBjfF1sEkeuhOcLTsRZE2pydh1GgQMhdpQpDSy78HEN
U8r/JQrz5mZ+MUCinewfTLBKzO+ertNfGqTjPf8kMH83XK7WCqpiX2zSPmKqxkPk
ky+kyxFPnqWMFFQY6EKHvZ761YUfxxjZ/i2U3D5LEhBSJ/leQ0uGXJ4qwyaf7hY2
cCONHQBbeR3FJTrHdw0uW+Pehnj6oRktkk60xoJLEpR1X5LkyG2sHfbqVQiKuiLX
MeQ5em+Aeu4mPTP93ThtFALV03yV0gqDIP3BRK1U+mETtgjILKzc9NitdwVpWDjY
n0Nwkbd9jLRo9JRjalWPtIQU8dmewaoGzjyiQGyiQQJ/lTqZ7sgfeB8FhNuPCsTv
i2RWgmrRN+fXquTfk1/F3iySf8mwE0pVG0RyrejQ4w5Ku5FCHMKhWvjQuxdYTmwL
OjtcwAuBZEWMYI45etS0K1K0CrIqo2j+uMTN5kEwgD57bljnQL3GJ2YYhVu7S87S
h7uF6c5/sJTTZH6iRTgsCqo4KHMVTsTRJsJ0lxYK4sUvF6mSVBK8hGO1jjHK478L
tnV7r/Ie+zT8Q2dVFSuur2daqOfDCixCSZoxheP1PCRMc8s6GHliaeOO1/fo0lZg
Gzo0TisCZs89HZna8Lb8LjSq3yGwdvji4vHZMw3HbvhTghlEMeCnkzYhXihaqCUe
BNS5whHe0edoL4yZRgj1RlLfjSImIOJ228A08f5WvgIMesNEG1wNtmaVX6FKCSSb
vCUZeHEJNkoP/BCLa9z1gWyLCzpy5TO0WvE61zy4FmBJlKNtuhfObgyWHmZUhf/6
5gxnB8DsJFFpXZYfwcyKPnGejjMC/JEoseXvwj8CtbLZWxybODEqWHecxe+K8imW
/UCXy4sPtC4Q124Ne/w2HC1cas+5rxrcsdLi5M4Ltsnz6mSTDpFUSjnhxuKC2fYK
zsXr44Bvn3E76uwwn38h0nfm7t7fl16Yb60SlG0D1xVR/h7trJVnM1L1CUi5ga4C
jJO2L5FmueG3dkxzZNg+m0RxaBqCHpUQnXsksjP6sIjNMzcfNEVaXfYNAtuTDxRN
STWLvdfHhKnBsz75rYU3xOVeMvjcim4wb8jPBzeXYhpIACWxihSd7tcQIzwDdcQV
N1vHtsKHEm8XPmNzSXTLgtse9FyPOwBPh/xohbNS3nUuqhrGT1dI02pEUH8DZycJ
WwQdwTIIi+mbyBrvJakmrSiK6fjUw0qyTuieeJ5lPCLt3uFZ77O/HAUofhV4ozUE
vUh/VPkRY8aJIZUW/FoVQVFvbPQPn/wBE3oRuZxJ6s7dX0cgiZhaf6AtIlK9NWt+
0TMYLCphf0qjnpUylnJ4pniZ8Qz/dm2zq+pQzpGAm2Y4Jhd4H+bOrUnpOJKt9DYE
WrvlfWEV7aSq90k68hF2w0n1yM05sXVga9j0sadxtSguF5rrTKakfJ2M2xSKUpWc
BxXeulZ4bfYeuHBt7Zaq3ZFhQZp7zaKt3mCfBNZh0S8bInur4CLB2dHKEsPHYNqQ
zVAVyld5vEKwv/7ojedC1huQ4xdi1rt0Pi5EomvC6qM1CzC6jYopFoxEENMGIz4t
tzkhA66dPIWIym1Sh8zK3RjqXxyKIMTqWc640L10KnK2v0WJPhmUA+/G4DxdExHm
OCZNzs8HHiw9FhV8oKBvFkO3yxbPlzhYEk3HDp51kgT8LUfHK7VZC5iPojkUtzUt
C4dDJj/YAoT7ATrtgmits3TIGpzwp1BdhfO6sklPmgLQWvPyndrJkXsVGdBzZsJX
TBiuRHwpUJ41RSQQAPgqCjsauPtnuioN/Nwgx2xG7pDkh1EaHT66yaZxL2t8iY6d
MibckS/Z85qZQFgic6wsWfOyYb86H/nQryA64GhWyN6kDqt0WoFgCa3WlBRkBVSF
mTfy/UxIQMoNIQJCcWLlbU9VvvNtDqPRdGj4HXB0KHWXey3ExMflSvrBTtjrhyTm
t2xhLGzzFdiI35+/+rwe6s2IhEuTKcmdcTBRhp7sRHn4eX1xCDOwG4L3/Hc/hIwr
odI01Q3dmEo+wYmvYBTEo5nuxnMmZQdGaquxVI+olWtsjP9R60tawPyqFRNVPFEY
QKorQQeIixrklBgRZ/z+rmOsSN1GqQmORFstN5fG6+9kzZ9ND8xMPZJ3l9B6BRXB
QbF9REQy3K+y/X1Mz0U/9veNpel8CBog907M8uNbkqdFHVFD2r3WFxUPxcg4oArw
e3yd342cFWSAFe1QaGCugpWXBMF8S1p4YfZRWo47DEbBehz3URgwW1gOSQiLCPGt
QXz7jba9imh3oQjIphSTJIVODBp1PIjdPRPkeDd+AdLUF1Pf3ddKPdhXaiTs4ue8
ddt9WhvY9bQjFfWBl7AwAe9gFOy9jmQueYUzwAfeu8YHNVGxmKmXZgZXLUetG/LW
GwqqGPThUm45Yf+6kJYLeITlK5WUwA3w7R2clOd8r+qHhjShdQkjZkmBy7CZ75vA
HuDE2eMph+2TdE0hfaULXZ20R6kS/kO+WsLjivcqleOk/INSLQES48gvsA2R76C7
rhYhQTjLJLFE9xpdBiWrTuv6rVnRHQqF3SBdbE35FMbh5WGX2ptgLtz1gJDg3txI
V8zeKUFNg6SytJz07+mz1mUSWh9WY51x1f40tvtlY08ItS6gsSw+kkS1DvD1uyhc
VPcPbRp690QcxPN8Dimm+JJcukptjU1jxiKmPoCq83GpQi1jVq0gCsBAt7QHWWo6
8a3Hrm+mI/Rz2ugxSPYt8CZYOcf/N/UaIjcj8ikrLRB62x2O024mhF3WxbFbyFsv
Di5ZLvUUY3DF0LWrigiaBL8hKBS3ZErzEvOa1pfbMWNnVjz7RR2rZnN4Cqqu1Rsk
Nr5OHblsKsVJbZQUYfv5aDDbBghXY/9UjkBWPczec8ijCogqgVpeAL5wN2EgRzv5
7oraid0kzGCfwSMWwJefd7Xjyo+7ThECDlRH147x2I+5jRDgFQHBLfZcDgsneI3y
6TnJB/k3Hyya2z93y8umkTPNB2RaZhXMEBzy3jC0cfOdzlJtfrnZ4uth6E7k74mS
g7BooXq46T5u7DNH27gSvGk/1DKyEmHzOZdgA44YN1WloflelrVXtwl7fGjEJ/bm
PEoebSCeSwD6f+uz3wVcnJqbZcwxVaPd5yw0InU6ZT7PzAL6Aqj3lkkvYLn5lkKl
SZZJExMHBKY8F+sKdpOER/zd4t2iycs/lNZ43tcILhZTptqhcl1QATrWHYHAg8fl
3Crub0IOK1BSBumku3BFsHI85dVfAqOwzVBSiCrFNVoLrE3ZI6sEN/PKZDLpC1M6
cZU0uMw4UeF9Ys84wpFUfngb030whzUt9HQl8f2bSXtzekimASSx5EMxIY3Wcil0
XcQjaHEUJ3j7fIRp2a5tLHCk5KX0Aj/h9daDH+HdR2D112WHP3U9WKB3RSilWApB
F+sxGdBlaIqHBzoKa1r9gpyc52hpR8gTp8p20qDTuOpw9cv9lunDyLLI+EIMOCwq
PO7r5qusVotTWVIVU0mrods9o1ueJbhfwBB3DckCaivfbN35coL61b0nCHddZMzv
KQegOfwSJNPj4St9qKdW+hmcr8v+LA6aHSOw8Y8XHnDEgzRMFo00JrXaq+46t7/0
NvceAAMpL57bcRg+s5FM0rIHYbS+0xDVQjMEEghaUJY79CI934hazVg7Im5Cxbu6
FjUdGJ5M5zn77tp1zXAULinwNcCQ0LRpTx6ajkOGQMUdud1wy2UG9LEqUbHQU1PI
jKVVz8sEAg17c6NH0PhFEPlzDlB3VxK8WmARjdva7L9FOY97oIjyerhBo5dRQVD6
VV77wsS+ingGMq4RB2/bHMfcS75/oAHwdyHC9XKi2ay5Jm+pQQ542+EelKXIOJPm
LF/jsWZ+ugrfjyTzJQiTXXNoOPhkikjljRhFer3hTAcmlFVvanbH6DvWnbMU0Tnn
kmWQ0soMa2T60ugJqcqD2NlaNubiq43OvvcCeFN6HR+t4RQsCxPLcuBcuwr63iTY
70imoqaF6lmOY/MP2dEUxrVa69EVzoW6a5LNsksabvO84jREVR9p1TkZWyuTMqpu
one/nt5xVPOUQ6Ubkc2wUwmoYzG2vxVlANpHrv5C3kw9bWNbiOQJTnsVYVUA48Bt
vReYsN81YRVNXuvuP4fEm8QuUIyz+IurU20BSn1A23c6pMbbL80ey0nQz+x9U2uT
BQKuEVHLLcIYynb8s6G+s6DFUytp+fCzpTpB/Mp3bKjf+vup6DieIZjzrjGKaonc
xR3LgAR+5ad7d79XLgYSUjfRgWTB4RvETsDzt13eUUmc0wyDq9WT7uMnlWd9KR8j
+OGfvo0kuGdQLRGf8ebKK92XwkOg3aCbOa874XatrAQyRtecupIgoxfaQ1hhpwCD
q/P38DN8Musl5AATFiuL60m1DY18SnePaYuFbrAgZRq+2NLpliHyuUxBRQNkaBWy
ndR5/yWdJklc61Fs4tCMnr/n6lLub5/ern8sMgUKADtNrXf2sLVLWJxuzHLdPR9J
HwiP5q+41isRUdXsp7oW/A07U6ExZ4t6mwnXrmOMws7/6Vgg3VZ4OgQ0ibGtcub6
C1+u+mbC8ou5sPPk3ORk0oHTDDYTbO9Xdxgldgh8caNlWmB8EIGC8zFXV9SeUFiX
J/steBKY/fA8g021tR3DFuz4qabKidsfgTHiIE3IHdygdMre6HFvFRf6Mc0Bgt2u
M7BxLgGWxipWKuUmLLzgcJYBkGZ4m3FDSHUoqQnVh17eI2SDAahqFC4ILf2LwLjs
HWYGpIivjveVe/ejslViXvG1IcokMV98Nu+6K9xBiJUCNmcgyey8LBoJbMgaLcP6
XSBRca8MuNTIPEYjGfWuGYi62U2923QnL1WByBSopK5C0olTfYSLAtQ441COpb7c
SZoHvo1Eb1ULAD1Vb4fP/KirBgT4zOeCDgBBRf9DKP+xp8Zg95cRw4HhB2UNgcL/
/eLx5uuiKM0YusMZtQs6QXmZzHGjExeYxkAJRhckbh4Nhk8gKj7GWtyGU7Vpz0wi
Dnai2Fp/EK2xdojQA5YMsLthBcfko80H2bD8u+R8AmrkBkCNGb/6M9Jl/gx997kg
WQts+vWDh0mhDEEpgJzFxfGkbrMbhXwl2M0OL80DtbDYVhDEKFi0lNjj+CBEsfZw
6bItu3amAoQ89MArYbdqh6jP5HWk9Pned8tBPgjq16aS+AzbfrZsa2LWVYppYVgu
Xs8dgZbHKYgcATNZymOb6UvEEzzxLcSnR05vPdjg8KTMMc4Af2n92mXM7r4T8L4L
vl+m4RAt1AoDzhGYO7NYqpoQ+uIR/HZp9Z3war5X+4YnnXk6q0SZp12t1Vc/JN5K
ImfjV5yrhe7R2jsano4j3NcWYEGhQ+8ZmxWyPKDss+gXjD3ArPng0T3S1G2KAaLF
N3zx9ql/wZJ0RvqZo+XYyHrhimaKv0dXEuQRPeNMuFLPB7UncrFXPaRHkyjEcdVu
cQ+YyeIyDEVmKCCCcCLm6RFqAnwNok1vNdoMT16tuHbNQbweZ6al4YUGV22xlV7X
Q/Lx28rswOAEV5jYh+Sux5xHui1sTW/AvBY+E8QTioV5sCiVAQTSE3O8B6F/nemZ
Tiaoc+zWwJ1RIUqq7SuK71xwo5UbvIngLkKerWJcQyx46MlgppxJCcPjt6Oc7lmD
itoA84okjzdPQOnb1goCYu4eRLUeUISvWRMO8aQ8b4FEftumYz+6lMApd6cZmROn
m05mtpKHx233180M37ICOC6UvC4J0Zo4aGYYEQKcuAPoS88znQDq2rzc89+/88pL
XcwcHkjZqfQLaLeXSu+b2IfQf+1iia6s4SpFSWYEZ4EM8oYjTHVma06F1C48i2F2
x8KuuR1grCG2e3U/w+d1uowUAplnwWciss6GO1Rz3QERisNuWoxTsuFONctiwm7T
05npIPxMFTtGP5Zi+uG1ZVyg9pW41pe8JvHBvkf9XbXmxjCe6Eb9fhF5m1Wno2Ou
djyjFfNMTTZ8aus7a+hwTBkieVJUZ7bm3yo9R8EjnOgi0kyH1ku5XSjZqM0DmoNT
w1oPD2cKnTnRS6QRX1poz1xrMkRCrJ2qNcWloGmNOzvI1c2lePzW+9tmJ0zKPGvF
qjLJ5c2ITkX6xLJ2GghbnnjgJ4j5lR5WL8RRTORYRE5u+qMxXLQhNovMTWoRc/bT
zo2VD78QXH2eyuquAiGITRte9WkjtVaWKk47pEE+YdT+PnRImRPVGpCZm+/KaTCA
2+97gmWhGAnzGWHbJM/cW1QNpqOWJYEwAY8dNNQTFpwfwkQTTvE4t1/x0OGDK/Yq
kNrVCvilmr+hpGkkxUIXhz0LHyidqmPs0MUZSB39f7GtV6R1e2ejRVesB44/YZ7E
JUn+tN3ylQVPaaYc3vN8KsgJ46udsG0u3jH9PaCVh5IrWvrP4+C+qTYm7ClBDDHB
iPr/7CgPwT3N3wb+k6+2oxw+ZhGIvotoqEIiRg4Q1Koj9RB0qJV6nv6mUB3gvCXG
OZEVjfHw4fgQNj/xJXPJM7y4uzwJvN1jND5SJ2R42X4tbmL743zj44KG/Oz1i68/
5RX+TnMlejYAri05irUg5fbQdRrSOM2LIIGAH37Gm4z7+k4SZdXlxEGRtwRbZlTJ
JOavSkE2pX4w2PIUIMVTi8Vu2F0h7Y0EDXp87PZjJIrdWrpkgdsWIrMk3/9PuGgJ
N99sG1YkzfPAhqi/ymKxvcE1EiwHOCf+BJHzZiBI7SSsesLdp5ZpTuQ8cDtnP5Ih
lwF7WEPhfWQOLD41pyDsBNe+vxJ/q8NfcMYPUM61blKdsSpwJxnHgD5GRTIjjGP3
XKBmYJGYysFo9OOJhxeNwbgvS5Ddh17tpQJVsgLZ2Pn+bCPvyt08WMZSmTPPGAUt
vvHsrJsZAbLOv3u1LpehE9QwzMrOKABslpVPaEMOUEU5nKeZLMvoqhJwW2rumkUy
rBRJMmPPmuHwMvnZzPo6z4kXQWTWHbxY/dZpm0v95FW1659Qy+xKd71hkiqdg7RW
52S3XfpCl2WV+LnxchH5gr9a9bcwReyxrGc0oZ9w2o1Ss8jtty2Y4c2Z/PcQ5OV1
CUz/KSup8YJn16ayS8L8vScpDsANSUAw/tbhMxNBf8RhxZejLFzt1ElVINXpq9T/
fsRYq8nSEQrlY7KTosccJN0Dcd/V4J/sfQS3gFFNsEqLvAA/x2m7IVIXPvs4tPuL
Fnzxwx3lXsTWDqnunJT3Tfd9NpmtYWKfLOh3Je2j1HfrGXUDOYemKFxhBUCBg8Lh
jPv6llTsnH0TJ/TO4Wi8EYR+I3aXneoX2m0rpDM7UA+y1Jdufzi3YPSFOx/xRHFO
w3Br5YvJ40R4R/lxRPIj09k1rb4ypAlWNwPHD0baNGl7s15RYvK5+ONjDjJz3IMS
f4cAdMHzWlhpgZFoX5ouocG385L264gTU1YMTs0jOMBwVqYsPpsZ5szOFLl0ZNHz
9lWvBy6UQ+QrK5uKlWXdj/39LF3rHV6qI+MgtTjyYJS1KAkOZgOgZPrft460nUgk
iojE2MangEwWfCBt0S4rzEhj+B/BJCiS0mz0MxBo66/UHeFV638bxj4xB9lrVp0O
PnMEQ0TzbyFJVrVGBMdLNw74vCLOBWg8UmS/8DaJ/DPoNDYjKU2NYqIXfd0bgR7G
f+5cfG4Z3y/zLV+NJs2sgIos8OMALXJLP5X+1lomFRBdrPSU8MFsbdz7QJFmnbvg
fmCXmxn3+Ssq7jlDk5X5wZ0NO5xjKkP/hNnVOwRS/pP3Y3kV6PmQAhDDJnD4DkwD
47J+rb65g/U9OB1zdFKOlN3snct5bNbtRKsVzqt/n7HyDOL5Pc4jm8bW9v6rYusy
DqIiy0eu/4g/OqnOa+l3zX+qZFIH3nlIcZ4hVQBwt3BowuBp3By6OexjxGVo7LpL
BN/pqzdBPYFOiG+Lv55mexzOJFEoAR9k9BlQlvhFS+78ZjSiWlgI9UNhledVatDE
ccLuSzLrRzujr7yr0Ebjs4l64wqkzIEWYIrAxZBOEao3UHj7Lmy5rd9scGmxhTHu
+Ae4twYAv2tOoVWotF94lbrrSMAWGJt2Wa8qAWDKF+ogH8rEzHgiD2TbBW/OMclx
ki/CffRlHaVIql3S4mBEr+zreVNTWeEqEtfiYKrfXtebBnNCLTVTT7M1xcqUfV7Q
SmGweANW3umeA4kjOw/Ag1NzeNADUx5xWcvWzr+oB6SUwsbLK6EmbHbPqtjmI3O8
+iCOD/wdmfM4JswhYcBSOAstbdyejQaNX29eHri2G/Q1HYu8KkSsgjlkD/f7i1HA
7nMRon5SvksZoTKnw8W4p8NGgw42KQ5EK8KlD+f3U/2qVEhy0gtYpJGCeacKbBJp
iyhVWjcWeWWCMqPh1/pAp5cgKaT444o9pQ3xlMKr8ifP56Y8xhG2zgxU1qfrxJIL
K3wCDwXCz/tHOweJSlyTXvoamfGFo+ocO6qhkL3TT9Xbbq/H5cDF93XW2LaA4we/
9Ql0/JlW1jxAB4i50mLcCQUuua2QhF4iOv8aqx3+qAh7JWSkKV8OIXPZPljv2nms
z1EVG96mkKK/GOL4+/5iB7gQHFUgrWqt5P9JavNr2onvG0F73yxZQH2lVcMjchRv
VsFWRMe9m1AY/wTttZCw6hYqh44FeZZmytvmoLRZzcy+zthItNOgHT8cKC2500qt
i44mj9FvMKHCDk01OZX/wvIaOHEyt9j5y7WwVOgEyw6AlsRXSZxnbOnwNHPdZItq
+1HGPWnYfgFvTI1npMGfN6Q9rv4HLNCpvo0MCcb5KmFbviKt3Zfj6itobE5NpK+X
duF41MiV6uAiTJp+jd15oRPexggCGbOADJC+LVHzojxdR2I53dl08d6lo4Vua1d9
yX1qobQnYr3aWHnSFhz6tLDhurq030BebyS58qSLlOi4dplZyq4a3GUSmocRqZTp
EUmJ45gOZkgkHKSuaDl4RryCaDAfVOtRrCMSu+L/m4nCyoGnyz1izl3FNE46z+IU
7INYi1jpvEY5OT9XEGBop/QEgvgcisiSajYOa0oRgxKRtHCIUbM2qI6dTkao1qpd
fHH13Di2qFbjK+3kVdrcgLUR7Q1YFZznLKVznl0SaMJKMW8mqrm5fwz9g/VZ57lp
wh92j1IHPaiYEIWjA+I8Nh6lrBnzpEKzhi+nllkMnDWU6wXnvsv1Tf66+/nsRLrT
ugvAdZeZHMluvRsfcIpVIyzA8iEQjx3EdRd/iOdayedSeqa4hGAtM+9mFqcKhUdm
ojy955PZZep1y9jRd8AWoXeQXx1C8a4yWYeARudRq1ysYD1/NWDcmB2IakpBqTBP
OSO0PUk6pl3Uj7nUC3apENsZyMGxC6659rZHwHCAN9tilJDslwtDDztKC5/7bniI
DHMJO1QL+S282CoKq3w++dW6zUpKv7rKypHkpeC5KQ7WMmECyX24nUx3IROdZhcq
KzvZ2bFOD1B2OiF2wME3oYoTDS7ojhRkbKT/8nN4A6sXJrEmCXwOxM6qyarvQZ+Y
7ZttOV/X0t6Sc8tcyIp2A+wuyhpDFu9EAJLpZwCCa5u9vHS7dUGpCFlCcGoLeXrH
/j4xWjF6NETMTT16vaggbBv7Pr0x6B+h9OJQ+dfhc5ovve+6WnzxhDXE+uoheHjd
ptMR0ySqPGn0KNerUKoRnJykQRoYE1INQrJPnwhGmengNsjvzhBd/IeRz2awYtS7
h78drR/zuiTRa5Lhy7wx3O6kvLA0AFzvQqh5oM1nwTq2+NHdgBUkX9dvfxGE3n9L
jLHb8j6jABUrByeNfiWL+ayWLOZCLOxxistJcIiYuzn4+bCxLTHf1PoSe3H6bPq6
7qnWoMGF3cAjFiInyTPj5zafSJNgbsoscgoc5Ouh8BYTLXnB6Fj1y/+zw2HEN5Uo
pc7iu8mCzOKsQwJXYjOfb/0zJrWXWtysLioKl2roHAM3ZlYtxVtBl1zhT+5CyNcx
6BSBQV80bal4FA4kLioU6mKlIKjPv8k7homi3RatwPP+Kiei++68ezhXKNyGa/yE
yiorIPnK4UVy8/e86tR6g4brHfxAtmz0OBX1g4JDQFruC8oFcYGKhraV/HkS7KBF
p2jfuiP7V2/sWPkqXYgzgfq7lWlLtDxzvKvOBscKX48/mkENNC07pYXUm0sUBchg
4fn+/Ntuk2B10NgXc2FexYDFLCa1duQgHgX/rApknxHfzgRsVZiPa9y7uDRBqy73
xDYjAhzgr2KXxsU4TGod//nWm/Pe5HseT7erJXtGtPAz4gAM7IFet4qaAM0j3PMI
QunAUwPGeiMKhFWWkHwlSBXcNDXGOvf2nxxyuGIh5ssvYL5MQhPChspf2TqAJ+GR
Vw10S2Hoq/z+pHXZfl8gMMt4fChbyAddO5VmESrYpbssKAlKr2cjrJQ82lFUrfdX
ry+GEaZ5ojdsGaMBGwMY3uhS0/vSMt0iuR/ThZc+pWMVgS0NGlcre2Uum1WC04TQ
zUxj0m0DSYlW0kWl+hP3IrDEL5fCix0inkHVyF0DIkqKfKGxg0uAaySZTP6BhoSh
U/U2veYWa6lqLEaI0SXL2Yy3gnHe85G7uL5Nr2U41rkNtVlUrRba2yIpy8y414GC
YTEHMibD3596I9uKLCelu1/0RcCnEo4u8l9x2jSD27i9VeJyGbVBcNVYgkkHt9J3
wtyEyDj/niTfhvfhziej8YrdlrmMii1wi5KR9/IPz8Tb+wWJodWWLJtS/ohnPHrP
B1iybYikkYsRTFTkYjdCuwcGUKRSPyz4IfMuC4zEXYt1WnBxHx6GGaBIO4n4wcoM
h8bmIHAGbZmhWuXJQ7afDKe+wltcrki1v1gDFqi+8aPy1DW5gYINqdGe2qI6U+ec
wiBBXtv66pvWb9nZFKowzD1oD1NeBFuLOyo8ifky4hA4v+Pn6uARRua1ILjBk4gT
q5Q48I0TyC/cXksnTdixZ+OGJ1pC0vGPb1qiHM+JUflAbSY8H4f4uiPjuOWr9c8q
zaUZ2p0r9Sq4HbvsqjAaKrkPSh1UekX0jpibxR+xpzUUBo4bh8zur5P/6z264CvA
lUNiTTOrSeJrL3E/RRGV8Z0+9xRUMIk4WIOOQYT+V+Tcv9sQ0NsoOxfxySW9W2IH
m0bz602+y7XBSEO5dbwsDnxaf1I4DEZVfO0tzfO20n2F3zkEFVgMkBrNISn0UVbK
rOstm0aV2s5S5Eob6qsBdaMSXZM6JM4XLtaDBWZxfYosvV4p//xaza9/X0gQTcyd
chFYe11kT5P0hmfM/zZ/4afE9SwqQDFL8110Yg5KoHAJkwG60eHGc1zgXCvEpdwx
t0kFCH0im9e4EppFSWm9QUzppskPFRKW/xoIAJlkYBTDtXFogeDJAKuu/B9I5hbi
+Y8QXmpHUIIaf/oLJoa+8sW3yx0dux5EKsJ02IkvQD32RZAiBNEQRfGrAcRg0svK
xW978Z4BSAyx19IiQ3wTFlh6WxWsyaVFF5xkBwNOwb0gXYkOtAvC7QbZVZioAToG
hG/FvEKLjOvlPgogdc7CSeodjS9CuTHRY5zdZGHzvKI1HTWFKcKdWQqqFdHTvODR
0pp+pHrWvNoQ6Ujmoi/64bfHlGlT3EW77o2tkfwmr0fCjyoHxYr7fLD4jY8SkFOj
I25JcsbZ0jsuDFt6qUOXbW8DmiXSyQw/nzoklaWqaPouAQrrRcVTMDsKcPorDKCB
2do8dNxvZRXrtXokEQ/o/jupUl9g0hJGybDZ8joW/lSUXzRAfdkZ3frRAcQ/zmM1
vBqtCUDGz4mJOCLZuqEy3E1LQotq3cyMUdy9eHRR0+qtcC9jcjLmJrBBjf+iLxp9
9qWwlmf/Q277Y/mPyFFt/7/26/7ZuSapIuFSKqbCymBRoaYXxvpR+/YRbPfagMHY
64witff1xDWuFtDPnN1v7w3rOQy+3V6+xsxPSrv6POSyCH1gjYc+GouZNQlKcsdB
fUfPo59H8fQHQGaAOa1gqscKVIrEuxCNLIhceG1bKOCSjB/p5SkVE85KMpSTDDnV
JU2HYT9tTN0pUx4/DCsL1bp2viLAZjYuLero4wJw71CbyNY4Zu6geQGJIBbycYW7
XFNwN1j3gqtHMIdKUysWtKPM7JPS5Gl9LCBmNTX/fwXwuCeHz1eEKC7OafRD/HrW
BiNikWZtm/GogCd6i96Kg80EEBY/kiV9klLC3eRfkHTOG5Z9l+l3BJDyn2H5Cuf+
YShnLJxf84P27EbWhOAr+D2oSrU4KvDJ6aBq5Qc55DHAyoYoQQ5lHrxCDA5a5waa
O80vMHYspU3UDWMKBLcI6WG2lp7k7a79nkNBbguy9Jtoqd925bgWN13PhYDt9NsD
zCQKtv7mWLHIey35zo3uasF8+Epc4RkC5fXWJdm8s2qqgOu1Iz4u3m6KzWHjhzLt
i+KD4jJjcYDaTNMhJrNa1+kMiNAhaeIJiym2M4WOta2Lq7tI7ba/NC5Yv1vSu2ED
DrIH1pZ5cYp4dusAPvANn4vq6wROHcoCVRTVjYzbABn4K/+2ffay3ac2v1KmlH2H
wUVCnP2wocgtTedbC0Hh6TzXSZOiBeqCF7CPp+beG3pz3eyZUHiyJSev6qjnceVH
HPc3yA5PIG3SRjih99c3qyBZOoIf+YzRfLcHiecfqjbqlEaJUprwNzFeO4xzgZSJ
MhrMe5CE/ygdcJsMKXinVahGMu+KRyhSsvjm2EH7+v4tkpqd3N6PwNg96d3YSd86
ccUeSkihGBnwjZrqYU+550uFCfAAnWl4rWvr4J2MnycSb55KcMh3C44ftdqoCrY9
L8vgwn/Inf8pzehA12yB8xYc4CrTfCkxGUJylH863Vo0oFuuVZNa2BWSr2Bm1dQZ
za6JqRE1AVABsU+mfYxzjJKck57wrpihYY0G379F8qtSdgvVZ/kHxzseVhJeCh9x
vNEWQ77WGa6hKOqRhLHt1dkiXg0zDdCXtSk9D8oNL7VzTBz6A1HkQPCcmopWZ+6a
GXcsdlXh+obleZEUQ8IFRT4InGJNaPOzwcf1tqnU2Pf2Us2SWHrSpy1jf+6uJv7K
zSC1zwwJWFlYPdnsS35bk1aBVb05CPlkLJbbvE/yfLurvs1GQR+RRciYbJRgO2aO
aAdoo4RZev2+Q3CDPYMfcSwaS3GVFxoA7QByJMuAbf14TOgc5Fb9yLDbT4hL8aTR
eNkJnC4adh+QRLh7B0k0557vIpyVkevW0LDv2uMcCU+PsCWJYVvo8sg5N+xUB09p
Ez8AHHBUk4VJ9Bw1kJAxdTMfwsHmeofTMtf+OMTcVKdoq2ZeQdo7fGCdJ1n+m8oj
wwYcKRsZk+S749Z/hjMz1N+z3IQYMRmqzoJT1NBuW0yx/uzndZWGDt0Wkudw9Iy3
PE2zXRN12HpAJVtEXRvo3ionQQOu07O6zyXh5dnFDuLq2I8C9S8fco9riQIPiufv
eKNIliaHlnxTjujH7rzPTqdPmYOndZVDMwclQ7TqU13vU+NB/2cOaED4UmXxt2XJ
B7ngpwxwq0bpTQ9inrA6+CDvzlz/XJWHGwOzhS9jBAl8VTq+0Uwm3q14pm5u/sc1
CfZqc2yF92449+IU7RHHTtUxsNx7zACeY5Vj2FM3iEAYzGnlS1k2z+qTyvgZ0kPE
qqe5FY4KvaQ7JRgTU95l5RkKH1KHns+LLCzqle8i3jbB8aIo4EqtA0XXxJkHYi1R
zLBdUBUO1AAKB6yObokPHGn8uXXcRAC2XjgbtTmKO1hSEfw4O1VcN/F3Ak3fKDl0
IEmL9wAvUt2tgn36+pjDsM6u95xRPYqmoaVYbkkwLJDFXHWVry7dkRwCaka5I4Qu
yFv7HG9XXBZWFGqYORQ+oJnYjo/pz32DudyWbIrJIZ/+vznceZJ4jD7YmkT3Gxup
m4U2jZToQ4W8V1ZumsahQ+vUhwm0A+Sd5Ktb3iqlYX/+3ovjNsGLvWtW5Cg2RwPc
ETnz5edvaif/ChSxUAxfq+wvN9ZGDno7to6nmbjcf451TYbQpZsiQ/DFegYGqZba
GfGlhL6XhQgeCt37bUgueXwKOvnYX8Kn9ByNGjx3SKlZvKxaGDslSUAxGizs7AUh
ZTrdaHkNtcpnZ9dGN1pPilmCZhjzMu5ACsZ9Bg7r54n1MbeKVk/KTxwwIpFIB+01
/kDBb2tZaffzsEhHza+QMvWwB5dy+MIElAISB/shYfXYoRpad7gm19BPowTZUSI0
KtMZ6LVT5g5fQp3d6Rpjbc3HddQublZ7o/EIwbMw4+ebyFBAkQFqeZHWMV3KuGaS
CXN6Cri92zduXQP0xh9iYCBuUEz/Ll7lfltDABfqJoBLMT8YcmMsniTfeHRAU3TJ
zeSD3nbP7gUPDECkVRBURYElOkYHBINeQhTpokX5f7KnxVYy1irnk/qwSmgZR3Tk
v9AEEWYcK1kT1yxyrqhA8mNlhof6fh5DoKM3jyI87oIf5FDhTO919YbfDVnorWNb
nWU61yJX9o9JqSTSKXYvx4weCEMHdkUmp43YtXl53Aoc0SgdsOssjDkUi98fdWUM
Xai59UIFrp/o8OOZyRJLIChbbUK7UrF9WY/kNKWYugXv/FNhXTqkTQQIOcqiKZgj
MMjJJ1glFf479fnHouPxbV7QHITcOkcHr9HNZay51dRGPVOzhtWVg6Znw89tv1Rn
HsdM3qgMmDnTInJFCFJlwYRojuKlToup1pIm+Q4/FH6/kqMgWbpy2CQZjsu1VJk3
9NJ9TuQjJ9OKaPn2QqLg+Rg/GJz52p2KdcIHqIn00+dxsNGcyUPltY3apbPI25MA
66zhpgMlKWWvBUp6Y1ru192Q4mrEDLT8ePZQhJ225iLrxQ2eOZi4gQD04ZdsAgfs
jzJ54b2GB/PMaXoGJgmvf8xfDiK/mLEAtC0bI6JDep2ylbge3ch85ThR3rDRz/59
+pSyyHRnMbMS3eRpnDly+givLkbTLlOKE8k0Zkt7YVSydYBO5Ao46+1QHH20cLPq
CdLaneO4+APN1VeoabSkgvp2SwEhlvWZYSCOnmtPVvUk+NvnwFQvH0nHVTLuE6Jx
hgbv4DjYmkqSDo5OQjRArFUdm+F6vNvW5HQ52KI3exVPEeT+B6NIHKTO6MZaqV4e
88Z3x1ZApP7lgXcHsQOnWzLGM6zQMHYa+9VxoJU7WwvVXdjIVsvO5RSzuT25X4TG
QJIbQYkDn2xNWf19TXflKbTv8LWvwBFZpo0zAjSbRsGHJvTpTXlHmOEjO0lx1GI1
TPL36rIGXVlbcwbPmClXgBmRFhAcs5zW2FG/s57Kkf0dECtteoNWJXXEq1meffxR
VbstVgSYbZNApdTflmEU1bESSNjFIV5Ff2iAIKAIoccoGGX068si1wXE7rdpeswl
AevD29WVtkX1BvjlqmRMhWjshtfXyjSBmAHMOM58OS1JVuYWXMVJ4qLAF/hqvjrj
nobvF+naTGypF8x2gp/USSi4wfsdMwTvWS7tACTQKQXHCzjnt/rEWAzPAdB/VcZF
f+xszPZ5lxe7CpQyMGvCuSrRDcDA44waRzXyWSwc9M3v9wHBzDE/lXO9qFROGvul
9lZAtE5u2f526MS2Ke4eWH7jrx9Fph/DAhuu2wAzR4541QjZtPE5erFGtqw8H0qC
+8+ZfHKLbjLWvgBIDeEgx2gIXFstQeQs2l7Y2mJkhaSGb7WMpiK76zHB+kXSzDxW
JzMj0AOwFG+RYSuwVoaWKtLN8bHQim7Ihy8P/d74BxkWiEO+wpywB5tJV22OTJb4
hsuqvVhWvo8C22x4tK9cykZF1GOxuvIjpmYVdUDqQAzSlyY6/Y0gWodjDRQe1T4m
9IHMhe7PVi1ABoCWV/oyFBjwxCXeKlv3BnoZwAl19hJ/QSZfNT6w4cXB8+venDRe
SwOBzCgIw3l+SaMq4G28e2DZBzRVPTCVI2f8ugasPiPhMFZzOYQ4E2fEjG7He5xG
U9PFC3o08sMdLUJ0iUpNixp8aGoCkWNke4NQu1B8E+Z9SnD3GoEmgjtIZhrf5Tma
P/05ozH0E08CUj8v0IjkOAa2Mww2/Yu0rtcp3W8aokfn9uXC9ghHVjySigyGOt4O
BzW2P/uHXI0k4lJn8ObESpmeZyJLRK2ebJY6TB6z4DMjSwXynvlyyHTfKs++grm8
agDuFBjs9ThIeagDN5L750/0iyvf/pg3F13IMVsCmYki5JnZpU1esU6uu/eEj0O+
VpjQ7K+qrsmfPo5fNVg/XG5ZHC/QObtGeOK/kbVCG7Gsr0e/XxhZEUN0bOvzKnd+
E/xtJ5okKAFxCgbyemq4BKFHp6CrQfxCLH2bi+SLfW1AIejT/2EdFdmUNU1G4/tZ
lSujYBv7lsnhHpFRaumWhOCE9P5rHGp8Ior1kDmDlcbdioXHiW5cZlbDYGVcd5TR
EHlNlVQ224FtioJLF3m8ciMDZ5/TiQNpHfeRryCQiLfWhM1jgwhZ3blOUb6qEPKO
8Ja78Llhgp4ku5sycXpeO72Xo18F2ap2ATH/kL6M5+Frz9a05myFWZDp+rCWdNFq
Y/mCiSaL9aQfkdX1jPLIqmaIj3eNsNI7RCCTlv+WegvwsiuDX2U/CBEK4ePZ6+fl
wVMt70LFOOBYgmWmZsHG7B+RfeomGTeIhlYLKvbu0pc8ZRSAu3bHvnv7q9KGpm58
hn1H0RCk05EAqLN9He1DcoyrFe/4v9W704C92qpVTKP3fRSzMisI9l7lWWk9eGfr
M4bizl4+ITI98pih/TlZB5BaeH6KPsyCFG7Pr2mIb0i4IIq0huaGJ/d/cBOC+H6h
80DnPdcEOLK4l1L6skzsn70RXofy2IdseRFmzOuETgF8fRhUqFPPCy+Z/YFv+M2U
l7JkXxl3RGFW+XJYnDc69+Ho/vezKxmqkWiI5+FUwNjhLvN4OwbegU0aqMwpyizC
viwiCn57hgV6jaVGzQTWZYA63lt+M3GaJsnIwdpcYDjFN90JmcYG8KO6uTKIIIDp
0vM+N9ZKQcGTw9hmM4KOx+xZn3V1aO8QAhXa3hJLzsLzRm0QQG7TADK43GnuOHnm
ACtiSB3/0gE+eRRD0ziN8o/Xi0B7OGq9P6JAFzVzOPNVQ58r2YfZIa+MDbVMeo5u
frlX8BCgrruZO7Gu3bIJaluNHl9ByzZxNKx4EvT0h2LJqlfCH0dqrkmZPMiUSJLd
sql5EhSobjDpG9rb9K9D6QnLyTBO0d2Jk2KWGpDdFyxF9XwBswixlZ11zvkFgXX/
Cea/FxI8bVzFv9haJuFzlR3RZ2bOq+vfvhQ0AG9tm8LGxSqAa2+lcbvfU8DI5I5i
1NymTAl3lH0lvVuS0qdH0hhWxAOTzIX2orcBpVjjkghH1Fch689Rsxn5Wi/HOgT1
iNzgigIveez4d9xMYO174O0XntQgeIdWmhfWF3/io74+NLJU2aiEPu+ul4M8Hr8U
kbK7bTLEvQun5Jfe5wGcbD6dZ/A0mIeydsa2szFwgx++74VfGR3I9V5YpaQGO9uP
98OaixC2FJGe+kZXKj/sTpmNomO9i1HcpG+STKdptgaCgzH98sDp/gr9izAtLwhz
geEECoPhso6TRWNgvympHeQ4XuFiMqJGch2dso7H5DdZ6YyQJhMqUdie2PE+QoMI
uE6Mzx0ZjDxs9qSmDJ0lxYclTAKV8c8dwGb/BN0tsFck78y8JwZAfPNQUfGO8AaX
UuheCEiYTz1b6lsbR7rRDy+fklMah/8ATTMTRLVgXwrZnMan6zjSnqKRKxDLVSy5
/RG0QL0hYYfYFjzceE3YH97tAzWZWIJqDBuROlrYu1utqoOwiWDqG63tar+i2k/z
Q7l5yEnQcCXGlpK02BS7hhm+DZGYph+j5HNlWGnTarHmd/VsADfSuwX8hvaPlbCi
JtaDeXKaILvqnoCENVFQn+GbQGeVAIyByaSj2kbxaIVzLnPVgH8glmLsWImCb/ck
JjxbZnQpS3c1sXLTJrrdQO4i4EEFH3vM0fYynSUZhVHtllwTR46QMbZLxFOndHNW
T/mk3ovVM2hB2O24wqWQOcv9njRTx1912McQWc66duaAzOn7TLqk9/JThQQZOI0X
3xEx9ywLcvNrLAWgLgmQMCIFM6/FmSOQ5BjcLh4HT1/vcb9onglb1XyWrG/9D/eC
Q9gZc4MerkPjh7ZiwBwO6Q5dcg/ZmdpUzslE+0pegosho5UEW8xiatEnxE9bhgSj
vFh9hGFuIfe0lrDVvzlO4kq+T0YL3OB6CHC0w5l1A6k9LM+Ms4DKPbAZ6XVSz2ue
StP/dxsQclYaJ2j+VhYwOR16sUyJI3FSyTfhpJUF0UpSSwbwTJYiICPKg4Sx0Vkq
HifN3FTHlyRh3h3eg9S2fLnOPZ4N9GlKPnopMwidNbv3vJ/hmMQf6SL0nuoUKJdA
cyXj19Owku1QSjQatsbUn92DDxCAWOjR9mZGl56mm++QG4nXt9gtynfEXWtKOU+Q
X5aM9bFWfJJ91G4qbzn7rjiYNa+edf1QxGDzSxchIi5j4WVMEQnRGCpP0d0J48C3
c1mIMHnzWx4BMf385ogNX7DZ5SHFL1LsBaYANSFD26hrlfCP6oU9gBPjM7f4EmF9
ZuPFHdmUk9g81HaJYrAd4Qf5u6N9wMa23CDbbfSdAOtBmQYrI4vNziPmR7Uxo7Do
LM8v86pmYGbmCeb/1ef/PpbFGG5Bk6aT7+/ugyA1QbIKYqXR8HabuiCUjBqUTy++
ah5b87g6ACOvWHCzyZ8YhVbUM66JUNtS1FvI/IqakAuLjf7w8BoH0HF8L82y88Ll
fWYYtKQ6PQpRttctYwo8kHanryncQdxNzDrlCK18TwgfN9V9L58kaYnpfg1a0LtX
mj+fYFFVihpWf1RKTU9NkovC6nhM+XFm8gfsW/nlRhvAHXIeVW9RsMzhtTOq2HSw
njp/vOh6xgbUgWhYfN2qhcQA+YopzDd2RYbzKyroePsTnKfJaURKriCaUvE7K4IE
rCa6rQQNLFea5tFdSmvdP89v9LsRKmGqk42pwFFF2LD2NDgefTfxgG+Fe0X+c/KZ
5R4wxZJzErsh7d1zDaC+Ve2BCzCFReXh2hAZG4a9u8G8yTaEj8b80IXqDQReOeuy
sOxAcrWaPQqlTRpmfRkFtOZyR3W+0MjERDvDOezcuFkGtVR/gyp99JZQHuBgglRk
wNSmg62c0C26zzE8vwlsQ/hBqt4G/7LBjo5i6sJWfHHFUZp4mmyaW0CP4QTfvTMN
DmXWK9Kg3ou/6VcxFQ/0Zf0hEHM55BOEqQDPdRz83hct4IVOkNi/H+MSs9giyFzY
3C7BkDWSmbaV6pwONs9Qv5f81TB4vmOCscNul8Cvz8JM13Fy/9mViaoaQ5WhssVK
/VIe0+Fxb2LjfeR2YUOaO52wd9mtghePm7qP3a28we4C6dNQ2sTSlD8Q228+gDMN
WSEfQPjr3rN98xIiGcIrDyvn6Xna2fPyfpKGD9RUlJqPKlso3piFSjP2RCMEKdax
ru75Yhj3QRdnsC2BO2ksMD3G/czTMGNgfsbHQ/ty8SdrlNa4z0+8qPEyF5PKCfHM
Ek0Q1QFKD2qO0f2KiylspNTa6DyZYoyrsiaolVSb5ZzLSTXGW3Lh5OQaKZRWH3Pq
c+fPnvqHaemxAtw29saR/72YKFk6ghcoZ5uFQKVVbLSaQqrYYCI80SvLVlr79mkB
OwXAV93nVci6rP6NGfFwOmMgHP2FFpi6PvjHIPZ4ga//FP6YTxUDbtxz3GIfcSyN
xr46rZquKW3H6NplbdYUKshZByQJPwXZowkllA8ZFFoRXt7uRstvTXG4l6vrFb3o
zzyGS/mfqw6CG2PRbRK0C4+Sd7aFmpwGtp305Sgz/oZA0XoYakOcXz9xYReZnug/
uep5ETM6msafracN31nEdYkEfWKdmvyB29tWVuKi44VOtiCeWD5CRQlwtYRBNzJ4
cmAOuJNdYk1zVaKcIS/FIgVaErARPdfWqOHpVX9cqyl4FRJEgzuyahOoptFV/96x
HRuD+fsLQyePz6JF3NDhFXsV9ywe7ii0vJmeHxOwzTd7FWgWeb3FjFDc3TPcYlva
jM5VUyjyWRZQujLV9p30eAO2Ap2sCkGjRis6Wi7Qjjk5t0mM7pGOHfaB+e8IdvSr
2GVYQGWw0XG2iGu3e/MRAXeGVg1Vj5v3lFk8UuDMiqoxDHbV7nsacg3nC7yWu9VF
dCBbKmAn8R4mIUAP7sDgVGO1mA4mdaC4MJjEx/Mi5dyruIlrJ/JbFaxuR6pMROo4
4tft5kWLHm2PteB/UtIP8rqZs6LzoaBrHI0LCOmtTwoAO1IKoDeGJccOb89FVzm5
gZSwbFmRD+NxG/dRiQZ4IHzB3smH5c/u8qcDwupKlhB1s5mDMzARSLzZEQT8R2ju
0A53mDodzFvDuj3YyI3ntgs8iPZ0hx066xCBD6O8ITCNdc1ZEiyCr3fOTqQpeAm6
5Xx0xP0aKdEALHQOPSzU6f2c/3J54br1+nTRXYBZZQC+hEPXoqQBAc3TL1MHIXjg
+tULTqQQvrOczjYkjdzqlmaJd9UZNonwYXn/fNGDL/zxLIje3/X+RfNg0C5mr5IE
PAbKh2D52E/N/mYQu295JtCFWhLCyAMOG6bPar5h7wtWlE1f85TyxXDkYRSQjcCi
JxoId5p+7KZhMQKQr4HMcZmygiZg1Scfc9Du9UkY8RT1dcmWXd+tMXKeZ2PyJitL
IUp8kwd0cWtb777Cro6iAHiUyf1TdXkoEz4B0h10LSTr7ezaRxPaelQnt9oez1/2
rxykZZYoZW4HP7H7cX0O3AXxEhpZZ0SolyDbeLbS+NE3GBr6vxHdazVKN4Txl+Z1
K+VwgZhU2TcV9bJIo5RobSHo6XUz088j5K5j8okCg8c1GD7HXmG62MVeaqPpCqAJ
U3qpqFqsdtfibJd+rRo2XvGY3Qz/T8m04DsvKgOaGAWiGpfW5exJEqhkfD3+9oLN
qJkEozBlWW8SBcl3Fj2hjv7yA0Su2G0vA6iLlB2bmAWmSMmYjq3bPd7+qWaglToU
dFhb27q2p0Lxj8W+sIeCBV3rij2HfVB63M1w5nxKq1pOMbgLwhuT4XKOsDwp2hSB
BcwZOCIamqH1/LRHzLUbDEBd7q2FEY3Dfd6Zup0a28wnrIBpiOVIGws1Z6JqLUcK
QhzAKwOMEiNi4+LETI8ptXQx0Ru27jJbTzE3YITW6SHkk1Uwt/FNofNKZx+klsw1
XsoVhGS6SQjH4gWBnzv65hxoslyoloXOI2E2Lfepilwl+CsgJnic9f5dFZrrrSck
dvn2oTmxIL0nrpGPgK/igGPJah3ryUnIRYB7Bt+rwNQkw5U56540oAnL2+qQHXl+
0AeOxVMjtja+cySQ2bFnrPL1F3vfCABPQgd4H9NiwAjpzY0GKJvWhqauL6kCPQRa
1O5isvMgPjs8uP+zlm9ZSi2e9ZJTSvjp79xAI5p8rT81Ys/uxSTx8bEk+mFuSXSN
CenKZ3nC1CcI429kmGKRPr4wcWHyjFLy7euObQqkgXGbzw30lUmTcRaDZpeD3g6q
Jajs1Tj2muDlKp0ko89PvQyP9poW+I1jiQQa5ChuOkbPgy7OczvuVSjLRSpkTNLw
oPW4F9cww5/oMAHvmSpW0zmLKgoAQAf74taZJik5qlaJkc4Hie3WElow053tJ1m/
500zTyPBKkNuOIWEiHYOQ4lNF+XQw5gRutwAi8e/rFMGOg+oX9J5wOSkxTkLHkBU
ejB7T+yOA04MNrM5nLf64b5vQr+8bEYvlwn2R+1V9EUN50XHSEAS4ucQBc5DT26n
8k9GsQbZM0ztGnKcP1LOknMyMowBn9Zlv8adVg+xCyN+facbCL5Mj5QqiQgf5xr6
agY9+4qYRQ6os6MmYcZ/j0TWnP6Wz06rnMXALXZPzw1qkYNGNGyG8VFY/PssP/+N
ZMAFgmueqozHnuNJpfi4MrwelIkvreSwTyTKtNG2WLVoObBAkIRLlie3XGCUwPtU
7MLZZWLlFhiqDcUYscSuyMf+qqHS2qxiN9wHaWa8skZziT2eQmBAkImEaJuF5dLF
53qB/zDKjZAyKjxxozvNblDzi46LJrcNBZDphylEspknOTtUb82thV6X57PcFJNk
4WJdkI03M2Ie4AltT3SZlpg2beYwti1Qphm2pqsbG54u+G4CigpkIHEH9jpqDz1V
AS6xRtYfI9Ww3GqhZp5upTpAdFB84yPdffa8cJx9U+KcuMbwJsPUlQ8xU7WOuHmG
6TYoWEQIAfmmBBM+f3RMAR3Kt9bSvQDMfaTp+B6w/INtD/vEpRFfHLlem/4hxACP
NDOpqVKkjJwK+NLQkNIUmLiW+vTWkcxGn0AAwRIEvbT38LRjYyCV6wpthFe5aZwb
UT139LWy4Ms+daLalTGbqPgHv77JgKRbdMgI3+R76fs4a3XJ4PwmUf1/0dg2icie
nrPXXDEg1ONRmV28bG1Vs2WSl67e2ebdo7bdfnM3gYGhyF8GqSwO7y9PO8ToA8ED
wEggGbe8cKsAW2logIL6Yba0buYPschEkBz0uD/A0fwfR6kczucxw385KyZ+66Ak
tGqQDKpVZxIYhE8FJhFK1PyCl1l0ciMdBw9Db979t/9pI5RXsIRxVJTJJl0xTRWv
0SRWwqT2rZRiAxrHQpslEJLkIUH+TSfwKe4O44yEhRdlctu1Kj09Ok/HUgoe9QMS
7YzZ+Fv7M4t0wA2iHok/hFFlpgOJdkBZMI1KsGHDdhI+CmG+C9rr0USEClPSoH1x
Gd1PPVVtpfoyugcZFwFIcAXUMV8GvBQD7iqRdNI8qf0rg8vS/MEEXK78rLfpkVjh
IMEvttjN+WPlYS0IaASVvRM5ilbq1rAP5/VaBvL9yD3b79RtF9z0DRmNoA8g9ea4
g8kXTmk3CxBFvYpMu1ik8rp5WbEJajuNBEz5fjQGU03C+i2vySycFSc0TDIidXfZ
AYhXik78h8/7mvgx/O5WDbN3lKkrtVecbBy7Iwjr7F4qlLhog9kmkqLdWkYNIT2s
PyVf7+jRrfgEmOFRh8itiUaRre2YsnThHQQjcJcpht6wqT/hGXffPqUU1UL8XWd2
/ONBMaZLHC0cTymM/x7kFYK0F7Wch8oF2amCRtP4z38Y9xxrkVJCbZ+nTaLUrF1e
qLxG3q/HAzBuIGC9TBi4vO4Q6SDIczOp7LeZrcyczzWkH+o5/4ToHWl+YzYdWHzZ
/4EHkJKS8y0ThbKxPpFLok+j5gmr8bWNTm0O1J8lJNkY2/pRj8me8xzqIxmBdEmG
vxUlTqsSj9lwP+V3zE4OFiLoWzuXKkjyic9YKpi87O99b32vwaaWVqxze+i4BUlL
D3RiFLLkURjDZubGeITRjqeyBmWacjjb8kWnpkCBJdI4rTZwP7yUcXcs4CtTXos1
jHvy0NESvaXbzWUHddqwo70AyBOH3uwc42xIE7bJho79HWOT8u/soRyBhv4SIGVM
jSrhlWO+um05ULUySjNfuYUvuy1t+H4GFFKa2s9IwcbxUq3umqj9xJvngcMmqezu
BvuJhI9uFk237phIARfvXSlfHef21kDkXiqB0iXGJjrgJGnN3fSU0iTWsizzJ6eL
jZXAT+phCYdMlxhDw1+OeubBbXXq1EQeemGXeIITvCSCJs0/xi3p+6BKhqhdr0ZF
6+I2GS4qrXndYyB+z7CznQm4UBuI8Q5zJ2gsOlIELwG0P4WNKLfHJpTvC92EaN7X
qx/ttJUFJEvDJ/sk68jSc5GCvwAQ2yXO0/ftimD/Sfhr7IlNSMWLd9gFewyogdgs
MzsMJKgTHAwSvimmzxQDf8JBDmkzBbbLJ5laWg2djVi5KU/2/AWpHgaXECqgocWp
SRlpXAa9/yADuWfsRnBH1nT+uA5hp9ff6hgy3joebmxsd9GZRjsH1FFszi3p60Dl
wShg5ZWDq5u6UwTXPsjyA+XBhFvBrmm48Qf20f/HJXET0Te0Cb42bqJp6jS8LJRF
QnhULp1k+Jp6EAUpnfQAITION5pxBxPzMqQOXNEKrQPVQLH2k2z7ASpa8omlAR46
rX7Q4pojNR+3N1Tf1qqtBXK/ZgM6q/V9nVNKWd9oqWWu0V7OQHl+fwmwTeZeDJPG
sWhFuRo+uvgbUR4bbqmLljlEeeKoTNMfsMdkHVbJk4NSO8HD8oG3K+vEOoxGnwBm
w2qeWvgHeeVk5nO7RwL6wjKFVI9tfHwFnFDBjjVAloP63zXR5ZP1SAkF0R65iPHB
GyLTTELuoQFD6HX6c2jzAbSU29AiLpxcd2pUm+CRUcu3OYyV8tHJraytyZN+h1+m
7cUI7d5ESc3NgYs2MP2KOKbvv37aDdAhueoGjF1gLWzfyN1jdM+WeJmjI+zBvrhx
KJsoqI2AhN9DkMS26mIUMvz8La3kX0hoKFzHaHlg3DOoTixt3rBLada0sp3ZNmIq
xB6JeAN6clWUb+8nsAicBnrMukuNA6rwAJ8xYBPR/GYxPG+0rh0gn3wwrasTzl3C
nuxDKS7OeCswkdhcR91XEkE9MV+7y4a6GZfhMrUZ/BkSyP9XGxovfKBlaYz+l6OG
rm6LFfqSsOlvCxbEmYSlt4Cxm0pluNO0FcUvW9+pUOYJ4pjukF8miQfCTKnym0z5
HA9mxW1PSHYm63mHExFPM1Z9MQw8lNfpYp8SISnE9QLkFM2NQTaqndzl0dv8Kynk
CXPqnChwWR1AuQl+2Hs6XM56Sk6qrQhDYfwdUjd1SaFi0JQS6q6VV1YNvco1MStL
vgHGHhMrZ5OGohcfmtAL2O4K6daAHb2dxS6WTMnga2WSMuW1Tn8UQyeL7YsbXmX5
JW/l1PdocGYgF0NxkUSzqPq2IARcYJ5fFRlK2/z9M+fZJJagqSX9s0lD4/+aK+UU
i9XlgcwPggSGs/L5ds/eLzchLbBy3UZDUoBrrnT0vvNfRoKra8XAr/0oEzIx9nM2
VIGf/auP8ZSw+xsk+NJvuIyJsZO/w/I7+J8MTVdHzIe4eD1ya3Kref3KxjbXuJca
4H6D2Kh29oA5+2fkJkP8j97/iSJA9IfK93KN8PfnRijHqrL2Uo0aw4FVWJoRCIbw
AP9C5svlmjyKeO+no4HvaYsbPaDCKv5Vj5x5t+2yVgw0FFvWmhgoLlaYekDDJAyb
VpGS4D9b1r6GmnqTngtOc7AkqhFKUu/swUEY0BhYqu0TdXLKKPO6JPpaoejgzczO
oYh5za41ra15gyNLu3EqoYNZsWjN+2Q/k/YIGyDgPsgiZxyCD8Tnkbe6CMnTXXNN
1HqjoFn9uqgbTfUSGy51KhGE67ZO+t9lon4JkAlFOh7FynI4tJnvSdBrDUQvPIUx
CFZGIXMhbpKZTo0cghWWcgtH5GvtUQ5HVLFcAmShIzQERWSNt1LspAZ3B+RD5Md7
TSMncpXGasi0VL13D02Tp6ERv9v4EW37c8rMCwsbnB+3MDZXRWtORTCNrnOPNxVg
jVE5W5LgrpXueklxY53YGAZIbfGGpJOb4kxkrwG8b1mtNgkrRNwToqrFdtJxf4qX
SVSrC5o/jcivXT1925vDZ2kN7Il3p45JOkx6L0JCqLqoOJCvtRKvCYLwyphTRHjL
iTbi+1urAlzJpl7GEuJFW/aPD79IPLgghHkX7fU64k5+PRRnUM36S27vMLUw2EVV
qadJcfElqsMt3IU/0/GaWCszmHzknARhD/d0KE/U4+pehusPKnnN9wdc+xSy70/S
/fGxjV+Izkih/vxdJtckUEZhYOrKlB8KdbN6PPqHEhzIsWT6suQm7s7s8idpfUh9
u4SlOjUOpBzySx1SBik/gWzDJOvMnpGS03qGis/obARuQFtSAEPFaHOExEo13oZD
g/4IavuZ0lnYpgvfh2EyXI3iEJkxwnKDxmc4niPDPN+UaUN5mLO1OCIRviM456eY
T57JyroZCOAaq/JNcG+Ssdd8mhPDRlud/7P0AAPiWkmEmAv+O8sbciy9ghDr2JHx
PqBCleOeJlIV1T8JsYq3bWHxIuKGtHf6lpIHglGB133HJNDKPJML+KsG0qMjEHiF
t/ztrivywPW9NadJX5QKLQTCaq8H50Y4L8zieOqX76+Hqyx7ir4siOptRh2PHR7r
r4aTWfpzLKXS4SZ5/+fFAcKWKiPazOHZBgq4VLdWvllsPrvXTM+po6tE2Dh5qshe
wc1ir/SXrtGyViROC3dtYNhtdqTDSqd4lH0nJODXncaa9h2Ah++t0+R45Y2V5njd
2yhOqQGgLH/89PHncRS4pBX8/pX7k1GXY4rRbvnsYxbHUTjOFDsm1s/iFI+0i6kT
WX2YPbQ7DhB0L6cTQ0MRQ78MUrRCO8pghdN9jAjGKDgULHYiMjOvH7PSfZydlE2v
UgIoOd1kdDp9hMKuNqdOmRklMiyQca+KNOYLeH66JxS82ZMT4gjuM+L4PCSa1P0Y
EU5IdnVQ8FXnypHFNbfwOpSWGnreqUowXeNB3Yj/Hx0Caiy7CHxWUOCkNxYNBJiH
aCqPvd+eil5F6Yal94FOGBYCFuZTGhhvUZY1JlQkhVeyODVHRJUrczjVJqAvoS43
omyO3cXA+G2cEydp6mykNG8ZTkv2U4GiR9/nl5O0HV5MHFNqtC8hIM2qykZ13e2N
HgSgIrvE3gM7YtBEVBw8Bp7+dUXDsIjiD4KiZZOKirYlPMAa8SmZsyIHxCD+ACBx
Nazcu0fTd0atudW5h4fYhd9TUwQiJNoGy81Xj9RauFgtGzAf2N+FemKbqI2NzkOR
Jph+yPN0TlejJLybDRcPOqnynWxTXfrHCS/pAIwiRvKtIHayU9enqDSunfxIrLb/
kY3s15FwOS2Yqs3BM6ezoR6aQ6B4P8We2IcKfRifeTfMhwbNHlaX6pluJdyNcttH
4MtaaNkFRRImMoUeLR2qZrPb355Hlbz/HHIFAkigU9n2SHseIT0CzqDpJRn4e4Ct
guRpuNSITOsmEDeoYXoj+HwwDIIYl6kIyrdoQB4gzlteSgeBuOqabWDJMU9yl6E1
bM77jOkeEjFNz6M7Oide7ouOam29VNgFZsNdxV3j1zyVbkpXb0OvmEjFSVcAvqNn
fv7frEzbIumpSPQ/2Z+H6IoNG+KWusleoO2UkWn/RNuY/Qk2eRobVINx8F+FyYky
KWNEOgWwzBhl0reMAGbuP3oV+VybaeiSV75QOK39bbtLYBbutaby3I88Uiyn322h
KMyooTc5EhU9hzIaCqG8ZYDRGGiYEYpWZdX21cANaqNA0TFML9MREeFiQqjo/Lhn
85KP6f00l3yPTH1GfVuQupawi+D1DlWFJoYwYosdPDoqmBJjWmFyeFhDd37zv3wb
UhlnGjzSKHAGtfyTIyhXxJ7ODZkkeeVq/hRavNtTutoRRV7XfFCEDXb51y9LvnB5
bYZ3OcD2s6maLTUFN7LhKRGFLFZ7B4qznADCfLr5fj5xyZpZ1JBnWJ4udihGciX4
/bvU8VWU5mg0+5ICfcfidt4pyfTZzrRh+T7P0uxHnvclndmEnqrfdj7AxIctDuQk
esOHAOeh8YiM6q6eXLrTTN8Xh/q+LAQEYVIkN/fOw3krAPQjQk+b9ToFHdaGDeAc
7JHUTOjbkeIy9bsIYTseNVqRfsMOfeliIR0pPAgw8aVhMwTqGZkBKswBkH9daMoO
n/92N+g2Ge72BUxzVyyH53xZ1qcanf7OZfrDxJG+w04G46TwLqsVhCMJOc/RUuvT
Z0pWoSIRr+2TV2OGY6S4D+TAiVWAPX2kMYaktCUawEwWoXle3+o9ia1WKhLyjR1h
nGjvtP17btLsLGhqvhK+J1thEoMdRUUSviW2MCNqcb4PBJrsdcKqAjPSmgBbEfeC
Gk64jJpZA0aTMD7OIKYAXZJrrQOAMnt5s78iqwPYNKfKfg7SYJS+9xk+z1J49o7o
rnKoLi9RsJ1X7aYdvs+TZcpazGwc41CE2wwbGC9+QepuBf9CV2zLCc5H3DtBaZho
3d4SmBh4y7TzRiSY3xbY6W0pJVRQ77X8s+9slQUIY/A1DfITp/MlBuF632B5Xmob
ptj31LqL2jOSsrWAO3RedptjaalF6U0wePeRy/uK0E6Bvg8AB0mVj8vVhjvMocxp
Zo0TdxqMo7/1RJT0zdZtBP02UyCbpqT49hZ9uJFdwoUBoqMBH1jovbb8GNaah4V9
m9O8SXPHITMlKOrpjZPtDHnLc0WTW7R/7vp2gmUiMOSz7Wv4YsDWo3X9tQ33cfdE
E0eo5qd3hcKvrIMy35NwOLnwPHR9Ar/KPT5q0koo3S1bVgYsNSFdy2D8hYSVFCkz
HItxWVcokifhNq3sCheJpUbSNCzL8Igr05duNn8Pl0ty2Jz8TRY/frgDNEn2fm6h
ZjLxDa5K+jl7oH127A0LuWDKvPBDjwupJvlHVTV7wzxI7jfK5L4psoG4zhaAHOlS
5s26ByDheCUv3ou212H9bckoNKyUGNipvLVUBDpMlOyc4jdz9GNCZ4ehTy7E1Nb3
Q1UJICGfYqjm/jTt6+PndvCJXw4czaMV1gx59ic6qGkDfwIrfWF0Rq5xzf+/jDHL
7ZYYDCj+JbNPokYYnP7wqdnN0P4D3q4vEJJy98kfsJm32byp+80avBqFz3ekMjIB
phQuDfLF2UbZhirZPd6Cb7+qmdFnoRrSiWRE1Bk5haX5vZL+nCfkVFJ30wUlWzqP
tZ7v8SHXnRd/UGelHRTC6W3aPf4ZUvwpjkzA1cMLLiXUT5u+X29eAXCP41mBK7UF
7/MBwG3JgLhilPn/E7obJSCi03rO4R11Luwykcc9DxLtYOrkY47jphuRMexxzf37
aEB25ThhZP2ElpitOx82EYQ/4jmEALqooS4fnFEAkIAA8xtz3V5vtSV5LKZ2MW01
JqfJ17Ddon/1BjNJhkUeAyQ+LFAcVJcSxxPuK/VFDIzXAK4u2JU3wCpva9HxF/xB
hFuie5+tKmww/G2+KcVGagQProiRniTroElyAxHHO0TMpdghN/5aIs3UxlRuzuKg
Fi1DloCqCwSmWFeKnirHs/h+y0Ryp4kcc85l9SjbcgDrfR8PRVkBz65PxfNlbCYu
MYh7L+L+lIH+8KeQqQeHPpOwd78o0h73rCHp2oQbSQMus93CWE6w9kdr+slwk0P3
FFzykacAednLA5pL3CIVk0umVg9cuTPl4iENg/8/cvW0oQXkG06ksOtDRd8tt/sJ
rhDy+dY1PQ0OQbZ5qI6OAYF66KgLSRyuBqXU1KA5StMh//1DaUaO0d+WfXqUwvRM
hU/PqN9US4Y1AgL79oBOL78SOfqwC18NK/EkoHnpcnFxXQS09kwKqmSJK6ShDik0
2lParO6TCE9VvOBRTW9ypfQld95nZX+ytEspppbfwjrkKNMIgkZVdELPNghAsuly
EhB1LFM/5orR+7V4zjUeEgIkqTkXeQbtvVD5SS/fhJsicX/FCVbkEAQNsrDmVQNc
ipvFVkNC4jGykBn1WHGUi5+VVwV+VaoP/iXM0MP5P2d3bwa8ZiYY5TRH5pnTIniR
mrldIibRq4KKwydH5fMgu14eEljC7dx6qrEDcc8pioeXFPk3hpn2CZB95e3jOKZl
zwyjTTCEPjzj7GfZeowjeQ7j23s+sZbi56zhwLmZBJkFTL2L6e7lY8pNbQpY5nu6
e4eqqy2q82FxbTwvNKWo9VGBs+khhqH43enGGT3pfjd3NNv7Sw+yYOsLIz+G7nBa
OT37iKR9q4BfTYMQV0NfK+t3kwh+oEcT3V4Lda7XPaNtn36Pfnfbh19sgUIlGXN5
zkep67h70u0O/3a/orvmdlLMrkTJtCsVR30snIDbCQBQwERDeIgxnoW5WGLVibd3
RMaDorRKMU2u904TTRPWx1owc8FlGSpWg5ozfKaDNwvpbQvwE8xGcSOs5Lm1XloH
iBbSYb6jWlGakIQX/bgzLljjFwhodMDJm+iaxTJCc7hk8mf5+d1EfNfmn/EgGcEd
oilmT2RtbZaODd3Mpo3h903caTGRayKLnLsBqtN8zav4iYJBKetQIyN4G6mDXvoE
IH3cogwmxrLwpIjgjPULGxRp5QCwZdiZefX+5sBdng41WfWzuh74aCZddeOAbaxt
qQ8qRqzCzXKnfyM8G84jbfruwGLkJKUGsANuxwzIbowZiiKJ7ZR82BZiE08A4iqL
cRyKEUKMgijS8nb1VCRmOQAZQQYvJXuOFHHEmkR44eypYL14z9Y0cRuSWChkj1fH
mR6WCGMWNBvH3DxssluSOdkAfEKczVvgOGAdUxy3Sp80fO2jksaAP437aCecRVoG
LKmTHPM/YRp6JVn0Zwuvxsy8nlsm3MX+v9F+7QvczRd7n2pVnSc3Ra+C9w01i2dF
G1WJS3jXhFsl8srAf1y1O+LDT4b7Jdxxb6jYQVh096dgBVWOyvjkVzUJu13Ky12E
DKJYdiJXQttC3VdwWM1bCvt0Q2BVcDcZOLbAQ141fBrkI0dhXAFyQHUIkZ6UAzMK
n+U0NwFRDSMdxYIKh32FBG3a4P+T7DDFK7esbGqp9Wf+0OTtdTF/IiqiYW+d//1t
QSIxxsMqKn0Ci9mlGmDdr0EfYPEXfzmO+ZGn16lEr81G+VKS9ENA8VNGepx5Og28
SCrQTALexyi2RW4JdgFu8FfZ8YCLx2HasMNJRt5eCKLv3zNE5O3fNSdeDvEB2qKp
N5THUmg5ODG48AqMvAYC/Opun5JBKI5d2ENnjzHa1Ad3t2slwXVUSAWEqhCSdye2
zKecNHMeS5zuhzSbFa+3odSqE113X8v8Xld+Jm/ONmyV5lbJqIbHv8J2Xn3J2H2Y
eKDGRLb+DhcTm94JWLdVVfGRmRpTYZunZz1mMMJt1tB7JSRajXts2fXmS8XMy1dO
mA+Yr0e6Sly7OSlFDzzU/iP1V8FT1XVWEw6d9VZpdQaNV+zDlOh+Wiopx25nU2pn
HwIory2PTatizrFJIAe/qWaqfhzdrcM2/ut+4v7yuUJoRhweCQjEZ8pn2UfMDtaf
U6iLt7/2j9IKFfrG1hlE1aTvxvy4pLVXGF49H87XpUekRb/ZPlW6J8eCiOGTFksb
1r271No4MpyWr0FdpMj7+5rl5FoEPWGbWVsjR6LS3Se2fYWRE/7YjwSpAEQHE0Db
SMBd/qXJdgFZ/A8gXY/gbwhiFMSCBMhY69pDr6kcfHObw72xdpMmGCCSno9T111a
r08PqtPhvGKq7+dhXZBrqLCRGq8n5EdEqN0Uc9kpZ+0qDGT6DHY1iyzqV+ryU+30
F1Rv+PZBp6zZ5x9EA//k/zI3kQylzIEfIuX3AO2/1TK+n3KFdnI0GdCAjMKoG2hK
bwP4WoyljLfIm5jmoqeD4t7DBwNx0PV2lxxcZMGwMk1sLPuft54ZWAglgj67cKSr
us5FUpmeTzQXCqY7CC9YbRdZtxoRWfR63xLc814a4I26r87Hmo1hS99XL/RN28zA
PP83iqQSmWJqyFTsBE/yZPjJHIFKbB6lLpxQVJ1SGDphL0tXKrwNCrO8RTS3zds8
/Kut7grMCJIY6/aemGeDo7wH928SJPGdfvwLVKxaDkKdRJCegMCM6KPt23WU4hB9
boleAMveoP2IHyOAaUvigh9tqL8HpOwvLe5SN/dWdJLn1pZIR6A9onf3UCo61Yfs
FjXlCJW0JB9bWZJFI3n7eIDp1XFvWX1SpcSZnreaJkrKxNtfbxKPAvv3EqsUVWQK
JyuJ2cKvvX13jJ4160F+55Y3QzgvKXgQa6d73Niuj7ng/6bZ4MFQNgeYD8+nQSkI
DR9VmW5O1Fzo4mIWmzRROxWC/l+cvt/W9kDVEzKFJkdSmM/ODifGtdkDf17CWPLE
VQvPC9LiCaO6vImFGW/QGHaNjgmA840lRDN92Dq1zVgubhWsEKc10sOM1oSeLwpH
GPzeEFEOzKTjeLwO8b20PZKFQWRzT2bokgIqx/TQ2BhbbLrN2jKgI5mM1H9E/0Nq
93yPQNSEDdoxI3aPsXr7YF2/hLqN5bV4/Ew24F5kZsLzV6xUgKXy7lsKKSSxLW7m
9Ca9ob5wNTcBEVGhJLetMEieJtX2tIZEOL5zGLOK8Szuhru9W5kXFJWgLAQMxumO
ZG6+FohyR6KRpWeeUkX0qh2Qcx/965sVn78WpRedhaLTykSdpyDt9l8Jar+eJ6st
fcgvuDrdMHM7ag1eoH4X8clgEEAOAm9gEOvmcCv0t5dxWDr/AzI4BhzUX2IVWrbo
DQ2F3KBmFjtEy+2AmOqgtNlaSJ7+TaEwomaOvW+SK04i/RBxsVuovUjCIlR7HqaP
u8eXgV4o2hHQxdLTwYubOOVCfEWMtW+iwtb4HS1qCYS5JrQ+rwEHCy/wqjDIeFCK
HNh70SifCzqwlApDo3D6dxuw1zKruPDi3Go13EfwA4z0nbK6L8S3wvKWoc3xo2Qc
j+/IIV2mMUdE+g3HFNZeFBbzBz8u9l4/jbpTqvHF7HKhJtFFgELQqhtcVlEwwX8U
DSTWINYHkM2U217imkRIitU2Yc876ZwafPLAfifYFuL4hBiL4TFo25CfV2bVi+9L
VY/8fLFYagPsW57g9lT4esRrdgx6XEV7xlX3fm0FvwbUjmbiuXYH0ey59DicoQNo
nfhTdXzzTW9ZUbCIWlcMcyEWC9SfLKtpiIAI/C19ka28U231qSW782SPKKmPA1H/
P/8pMJuyFUg6B5JMjkw96qIh1jGO1JlH9SeIZFo96Yl7TEa8JI3Y5nVFl6bYXvBG
qpQD21gEXzmCf+UdzpGFCeD+9f2feDuw9GwcgaYjjuF18PD7CKYx3FSPpDWSd/Jx
IcEuM0t5+Gwa14GAyHXEzcgo6F+RipZMosFNMb72y0IsM/8rciUhFd9wByRMB5HZ
XRLVMkxdkVcjJDQbwQ0FhpPPCmdZq2faj5mBXm9rRcDgCzsCiowUNp8XELhUmPVW
fp/anYHCQazf2RmDz0kEGV376ifmdnoRitfPXZZp5DAWjQJLvQjdvpHGJ91zW1Fo
Nla5mVd0aBWTMj1X0ES4ibY4/Or8qiBNkkmJDzqZxCT2Oa05+VpF/x8e/52If0jx
nQb49MiaeSihktDk5sTumuYVHB4DxqAyOvqm2YGOeQsy69WvZOoC6xBxpYpWO9mr
xNeglHZg+c7wl37EWkA87lpahfClIG5z0X/Z6v0CCWkmew7YdVfcw8PQl9z4CZIN
`pragma protect end_protected
