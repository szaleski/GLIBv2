// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:49 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
tFZrQfQSy+lOt/NASdEZT+siIZQeBos0SYYkBTddWHeBi4HkzsrcGFLDEm7mziVd
gD+1Xo+lU7fEZ+TDVC9Lyq80RDrOLXJHDRQgQ3NB91tyXoSlPoHHTGLNoBIDlitz
vpCp/oT8gWZjjcarV3Z6vmI928vAivFDrmeMW2wwJq0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 13600)
nKogPZG4Wlr+4JpC5TUt5c8mN2bCirP3fBhyT4on1a+7B1VIMHCRWkE/CRpzgEOh
kQxHkNaTdoej9Fi5QTivdap25SPLElnDyoupSe+d/s6iK+V56wVq1PG+s5PZGD+C
BRfeRFtt7IE06BPZIy3rBloXx0ik1hcAiAllW1JIBiZdezU/J5mFazvGzTBzf8yZ
6z/WWs5KjphV1dOW7R5l7EUsoQfrnTJBa+tgc1I1mzVobCUbUW6ISsyDUPPH1JUQ
KQshO2OVDJ1bnFhU0DmbILXiBzYsuvImeBSuea1XA6pNJtNsFvttmX7Ac665IRG4
JbbBXU8ncQTLw+QwxVy+vuNzrSsbOKKYiXZGmrR0tGV0uUr/9m3IbFxidxE93iay
qbAWlReIWC0MNtPZdlkjEp7Lot+Ms2CBRPghaJ6NJNbACwnIzgkEL9zydLhsVDLU
9mPhfZEibWyJuM3xlEzRa1ig8OgtHzsDVR6g/zRtzp/4G3Iukry/JsXcLiJ/L2/T
Kg9ouHyxoGaxc6bMQKCoJJ2mh++/vuLnXBwqPV0N4JuFFYQaQUkEKqao4cP+EjEV
E9FC6WAAAq+Cex9MAwKShQ/8wC503al5SY4cv2dlHPuJ7Lgs0NpZvH3z/cXuEzGm
OofMIkvNPxjbcJEIkrDpdbkSsnH5Dm5JH8AHKNSgMA8N0YwQdt8taZDc6oBkk+xg
4r4KwBM04lzY7F1uBW6hxxKIKsAv57q78CtH3Gmuk+Us6StF5Wapln7CdwFd4gsK
o3HN9xt+e4uF4ikUYEc8+SmllsaGuDXki3Ep4vRoyXdCT+rqXjodlSybzx9rwf5v
lvQXb3MoIpD734J8YR6q1Qjyw0Pl/HFHT8gwedasNjW3fgXNbAkEYEztv6yiV6wY
8ziTa2CSPkCGSxQwwux1ZgrA5c0OrYbR9XvWkeawugp5OJXBZVAFSv5YqJShcFBb
4EiPFQtTEPLpsJEgHr8flzK+aQL1X8Gj0TQZHETSYaNq8E9IlAnVWomudz0A10QP
m/bJre1otDzTitoxdb84y/LqTavDrqR59UFYmIhXYy1lbkqL8moeiH8LgMgLcXEb
7mnzk+ddRECISniUyHQcLrKM6DVwowQh3bD2saNYwkXXk7WoYcaOyvsx9p8t/dLv
p1nmUWTPuFcqfHic7l1xmYyRc/1Wc2eNvvAqZFIAYQ8HtvYrEk+wk8CDac+JsW1J
Z2FMqz4nMSQQroqeUZuEtBELQECNQJhEaF7VQSNzNOPwvp83OTWikng8YH3TX6fz
tEvf1M4uCboI3bF+gmtpQdLBtEPFf1VPGgXH2Gr+030XNhikLoyef2n/vAEryfF2
r1oC02GX9NcdNhzGA9OMfKtbLPgW6gMD5CG/OUBtjgcBbFgtXLqD6Hah9i0A5jpg
BNNHrIL6N2RR7HqHiYgiV8CvJD+qClu+XRC3QqQYNknyXYZh3QYhEwnKZKnU+yhl
cze+B1PlKuHrijq24uuUdV/Zu8+k6eH/7OALxMDT5h+PlI1AXXxRPaz6Pc9dd/G5
1v4X4MMdui65KhLWSxIkn+vRqLy5xa/fg7uVKRLnO0Kbn0sCBXLG247hP1CapOnw
cVCAAKaa8opZVWKY4OAa3irnRlz4G+A3PCixVy2V0vjGRguYaVIKw+QUbSOhp/A0
lzZT7lMycvaExSZhwui0EauHqeRllkMU3PDk/ipY+S/HPy+YGGnbyU6g2yBFJJYc
BJAeQnAnPLg7LpbMSW2v4DpABArjX1E9ZNG3wTVsaZ6s9drM+kLdKvmfDNmUQFym
HT1REvZpD6whRBiBYbHfprb1uvHII4OmzFcbR5bjLGmx2NCJ+KI28u2ZdaKroSVv
z6r34VCCm5KPM1HiGyrSM8JcP5hj6QtfAvm2sNI4CMxEThJiz4Pk4PZlWwJBiGc3
i8TuWoPDl52KGehBtoeOJmdC7kGQoG0ix0aeU1H0KhA217Edc+hWyGxyHrZWirwL
e5oy4CdHTWzlUAQfXEwG4PtBFII7GB7t1B4aCWwtBt6TE/pA3JgBa+gbOxrJ/Q/K
T6CGj1WsdHTQUdYgHhhfsrUGdrKnhXtoVda7CBBTq1079EXi4PdQXkC0fMBzteV9
JY7lWkUFp3/shRvYe4q3PFF69G/bjeqYLlGHUkNfMd5absiI3CtnLQNL9n27bbTr
yeUPjqEN7WbqUDrdWIfzzrD4o3o2FAmcOaSTWNmGohNY8IltmyD1DskV3Y4XDX7A
zLoJlaLxCsYSx0dJ4S07D4Q/tlT7MFQBhFLVAIhQTAI5RP+r/eBd+IDGPoWwIvrH
RZUI66R3WK4B+gU805gbDmlHFdZFF7n9zGWVe+If2xFynf1U13vPeOvvQkK9Sq9c
h5Vd1/tyRTQobIgEb6vNXAF3AmnfrKcqelSJQkFcK/yU/hKfYS1zp4n6sENTOYgZ
y8tnLlnw3JHdHv1fd9F1zgOPq47FHT7KIbZAFCkLlOMIzJN4X7c6a3faYer/E8WO
X5bhdiO51AChOjy9YL+HzBH/LedWXa6e6SdFp1iP3iV3Jx46qsuPoaCPXh9+cHYS
deESC8r8TPcEZS10fHT/ZPAmly1/ftu/0+aiwPz2LcWCVj6AbNmzaOX/L3lpKrrV
JrRZ3k9QxCrYKJNB7IHa9avg3LeVh/9/4zqo9m9cpVg1orTq5asYDmQz3fBFNSOO
owVbx8/kMSVYceYQ4m5N48+795SK6dzt0WryEjmT9+AECGq4PC8oiqydDcAwhSxg
4pFcfKc1cvfpXoCaIbGPBccBYgipNHDzJv1pK4NACh74T1svRJpGgN6xGLANc63B
5x8IA+mQe/YrjwNoNDC5RZTmFc5mss3WjpKOSGcAl/mDLZWEXgfZCKYgMw9LUu5e
gPwNM7zJaSiNqZ87qt8tkiHQyjDQZkXc85u2eqybuC50Y3E/tAe/hwR68BFN9rMc
VJAya+3JddCrGBjTMrtE4oSK2Gv7Ag7p1tu6nGfnJcm+ENeBGR/wzS9SRQ1jgnYl
4m/J9rZI+KF3iq/MNXF8VbtA7iVKWcda3nvsY6qkM82IxUyH2SVeh6BuXaJ6DX/B
PARO8Fnw3BmeOjw5MBxKRXVTBRjz4NIipNLyzaVPMdjSrcq2g/RE2RxnMuk58XVl
XldqtQ7eGavbUx+/UsluBJi5MjbN7o1m9NlJQqN6Crl9G0olwVJwvUI/3MMNETJ3
6f7iVPYLdFN3dE8UC4yZdh9xPgBbzHSp1rNkdaA17wfftDrunPnrkHbj5eQJTaV7
sd2u4ywBNt7XmQyA6XOTUKVmxkZby671U5xpXbYWSXpPpdMkq2mw8Xuhs1luQu2G
WEoWRtMwVrltuop5iayTVgYqzypznsaf+N2G/m0npE/6AZg6x7iD5Wl5f9rtQyEj
krkYzbRtxcvT8J0j5ZaI6//0+rW6AiXmNdWdcjVZeKoeJAkohmaHXH1wQ5+euwzy
IhCl2dsA00oKuu9X4fs2Ui4yIQUDvBcdNgUQgLEgOJ5GBGdMMDuiGp+8UgqEA6sw
5Pi+yZui0JV7toZCHiv5TlUpdhnrNdGYMBb463iQVCiiJQgoc1yEF9Qt1mKQyWP2
MgsC8p2wGQEyzPLn94kxdO6Xiy0ChZagWnWs8tM2y6CkpvmNK2Ak7wu3oSCD8K7Y
+M8VtDD/2Za4KLdl2Do1nnsMYhmrhv+bHxcOtBSu+cGDVQSDgBQaHBSK3bHavynY
KphrUgl5z9feAaSMT8iYMQ8UckXy5/lO6qDvfBy30TKswf8wPhShVPXjxRAfeH7W
w1qpVxKDwSMbAhbQBkXTHJt87z8PBMQYIrGXqxAZMTPTLEaZ6nZZ8tFWc+rMlwTy
h3Etol7+bR3o6tLt0cI/07ZeO6tnDFX/hAIuP/M6lC3zCLraSL+RoTQgoH4MR8BE
tRNAl67ENX62OJlS/htP90S84klVXXCnhVuZ3aLaIGfe+d1UI/w6EgmMXHyYXL/a
21apNSHhrgFrZsvTBB+XDVy6X2pPfIGRJfzPag13zSL1zunBa8IeUfuSX8LDY3Wj
O1gYsKXrqTSVWjDctWlt0CLfg9s//BZ8RPrBvn6BUEbosPGHb9WY4Sj0g+ovzR+i
7gXxsHFKtpwr85FoLN/z7iUWGuJhpOhMvmjFhuDuWevwSa8ukNMYhsJqjYlRG8P/
iZxR6R16tCUBmEQ47hbiTGkofIvGIE0c8Fle9m1oyuifu2+b2M4LxvyuOZE07K5Z
SpX8WRclrS/Y73Va69OOTnuL1x/Hl0nYxLvKKpi+xrM/9iBZJoC681rhFQTeQEv8
FA25+67dOqra4/SCT9JMWpllJoucYccxJkF1qbbJ6v85MxGWg5SP/DYVtsxVY7hd
4ICYr/BTyiXnZUfdeKGSNMI621O6x+SeYZ3vIW8sIWamzOaJvYMBADPFNOz0kLQ/
pz3ZWISOHl3PzvXbiyvCk/U023G4vYkbZUayemjstc3+oJUHuSgqWglw6+WYfQ/Y
eBJQCQKIJfZE2jYnpHHUQKexK+6X4xqjIRztHGqvi5eW5Gc1zMNatNxKCUZ/X6qd
p72KEc/cyYhe+3hET9FsC659a+qDv4puaBi7Ig1dLomHPFptcIPilOp42UmNDH7M
9c3JL/D+BonKEdkomXCLkvu8ByguVkVwOpLy3VLIGQSZKAqND9Ed/DML+PT7tmL+
126uNGvur/SQctpGlORfy9K3MVPWUF6Tjhfo3xyUlz0SR9B/zH7P8rglJsfm4S1C
69tud1eSzLkSDAzf4oH8MD0NsYM3NUXG8zbrrIGzcEePaZkBev3qdgTQXFFrE/wS
WFWLj/fMUMN8REv0xRSDwv/RFLq8hEodKXfxEuaHUA35+Lx7CSW6JvSRBTrV6Wk2
LLj5UaHRtbXPKWUpRYfICcGr8PjtwG/FoksBYJtgRPibUm6Fk/IAtngr++9oUhZ1
/dqWDtQ2ns1HV947ecFiYujkiq1B5P96INYBwBRkhRoypyTSySL5JOPjH7KSn+cH
uGfj5Ze0QJum+J/60yn4hrapNsa9tw+h0+JWIFiuTZX47xpcj7mIgGKQqHJYnQV+
WHIjpNEc/t8vect5Pop9ocdntpvxzE4QeqeLBCZO8+OdVSjWN0SGrSGlw6VPVR5a
IEfGJ0/LexlMarN0O6u4+WrAJjrMBC0PEdpEgBAcA2qP/8I7sfenKBZr6c3f7ycu
umPmWDiuVEJAvYTDEroL5j4Z7UHrLx/jyIpCAH7RQKaPJYHeD/QMdqo68yf17l0h
I78OlFZOygDXKscBZHPnN55SSZP0ppO89X4t3Sye7Mgm3GlDpqQCaNGqgTqITEO1
rQJZhL+ZyboKTNVE6ompksNVvS7nFha/ah3hh3GKrMjPqATmocZelFozTETMMbO2
1z6J72Ytbkpp703eGwD1cnOrwEn8j96KDPWZCBITSAVK47eR7RcKNB5CYKak6Yiu
10LtkMUGIpYdS2XqoAMDSAuC1rQ77PreKnqX+kAIY05IRHSypongsM+/AASSk5eW
LNoWChhsmFa8B+uEtTj2QOWKgGi4u5o07lBeuYHZ/kC+QU//jdq/vZ5QnUOhZDex
jS4qrswUDZ09+yNWImqohKYs1FBso1wEuL5dyfd9NaG/8+evsKhkYj9HNmi8C/BK
do76acGSPYLUErBoQMZkacUGfyY2aTRKXy6xIADt5gEptQpPl+HtZZUgs8Bj4khs
Cd94IKYxSIdwgHpLK2jN2hLE0mRFioRaPyuAIQrS9n81Vq6i6vJ9w+0h46diIh6o
2ucvjLR3SpD+JO53oE+qlYftbGmhYZFociJjHnHE0iq+fTWZUdgEEgjBzAjc5aI/
ecXhZMLGiuNHMvnNxNpGEHpWY7Ujq2zNOVvxO61sIEYXHkCE/k2x8MrlyO6WUeoc
MQwH9dp66odpLcEdzvHjfzv3giAQmE3ADtln7d5SxnUk0F0+yTTbxXc2B7tcVM7I
WEoCr96YV86cnycg5FyQsXNQ4EomyGaY6TRPJ6bi8u2Jwo5P0zjCDcsv4oa3cW3P
IncDEaCxiMZ7myJQbDwJTr0EjnyCnnwGnNAwcU6zwcxndgcnx8BNUNvBWglixSw8
pU0YhI6AqPS0sOUR7j+WBuQVwz2n+cg+JLrmThPe5UZ+N1y5K9YKyik7H1gV/NTV
E4Ej8O6ZDDeHh5Z/o+49vtqftrC4K5Nae38c/xmezGnt9eL5yWI8F+9yhwATtux7
loD49TW45ywAFOYOfrlekh7lybr+V5QvuFTYGX9AviV2uwFoPmPXVgfpQQHcmV8d
9B/53JVGCBFwn5UG9ziwv4HZYzzXBgvp/ovETSISh9hXY3vpUkFqwTERV9c3Dr3s
v96WSqnh7GP+aMV8TkjCRXmntl0E20tKuTYxm7jia2ukfNnaNNa08AwMMPMDo7mf
OrETbpOHjCc4YNFMeU1NYt5BC9zmCC+fxzukhSjK9dpFuJnb8l/SLFls1+j15G7s
RGp9LcrzyyUcT6du/sEiKooBhw9tyZZq7GioTKNreiYjW9tViiB67W2tdMIcOsKc
gComLiTuoAsmJhyGUSUWqeI9w+Ouw3i2hU2Y/e5rNCm8PzrqnHhRga2+M/uEu6yT
uav4B4lY5kqeGLMnt5XG79baeoGrrBL/z5xlFwTyoT2FGMmZ1kN416W9H8UOdjOY
ZMb38ubvoc+8s6O0t2aJSQmWjqvKrrJdW56r2oMHb2jRrhgYQud/qJOdz4dAXHTI
FNRBHDhEgQC0qsUZ+EEZTCaYPlcQvRkzQpiKS2xenXc+/MVzxl1rY3SDxfViD2OM
yBUOpsfZFwtUAuZWJrqXF4lxiyebsdkC60vj3nkNAGS8SMH41jYNqLxR1kxvekIr
v8rLzxX3I2N3jdnA3/EM8U/zeNybxhRRDRDzxm8nzVo+CK2EmDoi7zwl6j6isQ8L
U3prf0L+qmJgJXleHHEsjySKlkiqN7Xyjq0Z9ls3jg1LPlRsEMPqxlYVplLRwX4y
AFHbyC4ODusvdxh7VN15ez+7wurwa5n1Znn+EkOm0/bwuoFUR3rxYxaUYhp7zR+D
5C5LdlBp4hwc42HbE9P/dKKJl3U6oNPg0X9UktSMm/rICOzkzzoh/SYThG0LA3eE
ugB0Rlfjvj7P1ZDOp8u+u6LtsX3FOHcc5k0+KM6X8WerQtYtms449zLiaxWzwFug
lToa9OUJ1OVWk49f+/wuMiwwC9Ege9EidfYzZo8fd98NLx6SmS7VEKPfPRXyMbWb
WNEQI8imRfi5u8wp7zYREeyw4MaNv+GrgqRQmqBejpFXg3Vnx0inj2EedZ7WQiLX
+yw2ARZt2+0IJW0zbnng4VFQyI/sS9n3dGaU2HotinXNzgDE79msRardpBXI20gJ
DMhOlCrvZ8NvUW2IxWqz37XFKOravJKNewj2aOAhOpCBtOZZsYZo2hNb3SxdFhQe
4+gYVOQf6M5qVolmW7aZaR0eg2K+ehW2NvGbtqlqv4WY9chIspaSBf+O0Cw4jqK+
rsr1g+iDPqfuAL5bMBZ1j+5z0nIGXFGvMB2WlsK1dS5GN3nAewbF/Ig0JoVy/TSN
Rps1C4OKGL1YmUF3+9ESQPvEYylTeVpl8l2t9MA+wD1uPKKCsDaJr8obwebR/eU7
RCgOUHcOaFKt73szThf9cp4ukqWZO8D9JPoa9YU841zd3E6jBsUm6oxN/7QWeL4l
bORJhRzBsSXQKRBY1C5tesoKLfHpt/I0aqPrrGbsfWHuZJ7S7dU3D59lmnkIeSgV
8Xo1+SUbpq9E2cWP2zHYLDbRjQjYzPB4PcdYcztafLxM9splh+6yv6xyV5FT2iec
nQvdfhByM6NX8VbGVjc0wA08oHlUoHdbXv04He9QptmS3AtvryXce0lSv3ozERvS
ZILU7gYAS2ruypUEaKSuqXKqroTi6J1RdmllKQhoFSDERPVL8PaTi6Jf75u8iJMW
5kuaI7nS73mRQNlqj+ClzqCjQ+G1AtYmL1OAYdBxVfKo63OJZyaHviLaUivQrAbD
Cri7VSsBGaKICw90V3Nqt+XKHzJvs0XNACyJiOeV5CdtkHto4BF9+kyrlGHlisL2
1RtXp9soK+yGqLqKyx81/i6lo5+HrNU89g/zLqnlz8ZP02w88xuwXkvaDnACl5em
h5uUJ3SMWOWUj4SRErkrZpGZoEwnTCYRxhO7buH6H+T3cHwjHenh2rmZABh+yYG5
IwKaiXSgAdKk6WFo94Chwotbof2x6KjHVlexlsu0KstqdlQXAGCqaA6IxG4MgOxg
pswQV3cFtC7d9YKW1mJT5fVIWA/Ts2iTlVtpRFKunursLJztgoptZoAyEB6ob2Ux
QlBJpCADMFR/Jdh5/45ZQHGoX/By59UjAaPQryPaqmK84j+SMR8r8Fbnx3UAQaJa
J7ofeT+mV+pPqr7ub7dPFRB5YvM5CBJEJfleiPj4fM12PV89P2NEeMm9a9S7WBwL
QtbkB6oN7St+xUu7InjxGAVak15KOENeAJ5z9IX9GnOTJpKX4PyP4HWPnjL5JAem
/eM41/9a+T0WWrs5jn4l6almCKclgSe/Vg16hZAN4y7JyS9Dk7a31mPp2P4tLKxE
DRpYO7imbWYj/y2hH0YJ6nIhTa8bLwppnpUmMu8o0hWmTXXsZ/T3Tt3A9dIDDh2A
DPjPWQ0kE7i0BBMui+8Q/iVY6UQT7zuHy7HPJjVRutKUXjFzv0LRZIJ/zy0nxwoC
t/gsjjqSkaI22MpqVD6A7U4TswBSYevjS3AFZf3MW27tlUYTTVQp6je8r7ubNRwB
8scIWCPnvaRf6ag+d1U3rQvF3aW8usWSx/GuUxsob0utI48DJJIFFzCl6SVNt2mK
Imy21PENeAnLoy7QAxFQTXZWRQ4dkLFp079yo05zuIar1rBH4p6JU2JXvEFaUpzJ
0XZt/3VrXlqlw+k9IU7V8J+IrlFnBgxwgN+gvR+GKzPGAJ1SpHDegKWGDV9IFxCf
3hhxgqTTDqVPewoCTMNOAG4QnTAePCVi6mcMZHbo7GrTja6fTmxqVWJ+AIXgEohy
AA1zyH/fhElHrXjKGPfjYhz7Wckf049HznPqHriTiiioW08pgmXoVFBO8jXVck3q
NOZ2+W7a0x6jvAkqQn+F0ZLxiWCUFhE9iL3nUUPo09B3/nnRCd+2PtZSQhKyPgnG
pmliBSH9dBsjSTA1J0AzXnxm+lHUc7+wk10rKfi5Dxkjt7z4YINMxZcWes22Glf/
rmjE/BadsgW2tKPtmUlNc92kNbdQ+Lbq1vQaV3lxlE3eYzEet9wML4YoDQszIXNE
DuALwSqFGnxzYl2ykftCZ97AKp6ukIFLAwFBFK6OtK5sp3e+Qj2haMzWCJudKg6G
UVcAmOjaaxXKtcTr9k0lKRgG2g203kz2x4j4f5/leOr6jvSs46ye8YRA5OK/d0+4
ZSbs/sEX6H1LEvSz3kRvd4zSSK8i6FhbIBgf/mVHNmNSEIYDSgDIgB1d9qNNx6h3
PJfBvmH0a4aiRVslKNIuDqkgcZ1BlMM5FXolhtZKB4xYe9n8KwiPY+q6HmOX60EI
nUw/zeJLa5HgAARHpZrWoQEK0f6EJRKbdxdhIu48kSwJT/uAsGBqsGQnoU4BDaup
yckkIp+hkjXVWKk8ZTxMWk5PZcAxJwdWr6bJBBV1FerHUdYa2l7xg8b7b1+IUy75
C/hT3S2r/ngArgHgwnJ5C70PJNTZRled7XmWh1P7xB9AdnZJa20ljJD7/jTPMJzo
n9m0Y3WeXteSafhQLMQ9WUDdalshucD3bptWPFu7L8yEg7K58xR4YV84LWO6LJYu
w4eG9nFwHrkHWtPjWRtLzZyP+8XseWwH09yD9U1giSpJEP+GJoH/QNglSJAiG8C0
u4P1WQd9qvSVlfFyFuLi3Ec9g1nXtnl8mHxWyOuIpfkz/8N5MXnT3MmfqYcxa8fD
pmC9hWC801uC1T3SjVYm/9SKibyRPG7Rkv633Txf1XNeAnlxOcsgV8sDoCJzyol5
c7y+2dx6Gtam30s6WhkjmQbKjl0JkC3+WOfJBi0qP7g4IBglqL17eVg57MpmdAi/
QrB0QxvHPEHV2HyqQ87QGgvrjbLzM4muqxUzCvQH5NAwkWO5nFrRw46Ot3iRvW8b
hSjP7DQw6RfBZLuFQQNOp4HmhpnhzycokkYjOaLWTvbPjct9C0eAH37/BJe1DxI9
Xr0x+sR/hhEhgMv4imfWskryhJT9clgTQuAx6zYE6crWkEARp2h2lOljxSD5RmJv
mUnwkttNU0AXOHOiPiJqMUyBfZv1owUqAqAxKzZCScJbbSq+5LIH7xLtddEqAi5l
85cshYV7CYnIMaFipC9KW4IHDBsNWpCN2PLNdpuEmVaYmpijfcjjkEfmoRyPqDa7
n2BBq/qoPnk2hu5MhgPo6xaJdw5uD+DP4F0PcCWSozsZpjb7h8Qf9d+SYkcuEsru
/OYouLoKg9RMKzm4vmAUy6gyUo9Cno8TTjnlK8mQOaFepxc9JMC5sum/So+IQ3Zy
HAnPPwQ2Sv31bYy8yLErQdX9jYxQbs+e3++Xjwo+E02RPQZdW66en+PfSXZSlI/+
75553a76xkVnaOz3oIOebBvkWg8VYaxx/eFeYDZT0wlO0j1BYoybjfKW0LmNPs6l
Hct+JN7QDq4ZeV6ZwJhhYUx/TLOhYJlybxVsS3zPSpEFrYYxPUUAwoAIxwBDjR2Q
QRtpenTyjxqN13bGEkdY4rJ/z8uwXcuC0fbqi/61abXC2txoFjSsgkMPvwZWG6nD
d3TmPMbHQ8TAddcj7nq7SQ2Qc+zGmAyMALL3Z8ctx1TgzHmo9vGLnvnzkH1Z73Oo
sDt1saYW8op7K+L6YUVQVH6fzdB2v0tSH45wwy396eORAyTzlUXcogJNgMLdsRKZ
PxZn5oEG7Hu3ILeY01YrboShetRAG48vpUdLxK1wo3313knYj/gtjDSX3RoPx67z
3YyrKyOk5C4Mh63nh6HAyFoZg6Uuf/DtHG0HSIEG1nE0OofEDPVQO8nClO3vx3Wg
bIbbPU6Qnh7hQAPbyy6Jn0ILsC4PLWU1eUJbEt+9ySYQJMrsx0wIKpXiiQVe2hSs
epmtHg1cxF3yTxKQJ7J86YpSjElS95fDj0DjeDouewftEWSYq4+ouiOQDj6LD+oc
733uarNVxRg+JbzJXDwrBEWihVVy2tALrS5wW78Obxtc+dBScrMU+gyKUO6nEwxz
7FgifHCPLwj4S4nJnBH9Bt3c+rA+/e3wdK+wwzbuTnFCEZ0KAdG+sVhPsUiy5VHM
gYEndNQ3iAlzHJfXqE8Ypb7WcdDs+880zy3s9vf99djOcIFOZdioI0XxV8Y2AIcn
MoK3s5ytdM2ded+gunVgP1DY553nNNPnaW/vRfm0v6l/oUuNmeea8dYe4riXh00n
4bfFZhJThYwTjUiwWdh25O8/A5ZZeG25ri7if4MW3cJLVpk8p8kox6jynjI1GD4i
AdvUZExsxdhs+vusqm2+TuT1M6F4V1sUavKMGdz077/TXci/TO+zHEq2GsGVm9tB
69/CMqaa/QjgIHDjL65YBpxBvfye8qH3d78tw/MNoEsIxpCjte0T/HZdkfR9Wl3k
M+gU65u0KuGuBrci2GOhr7QmjITf3jsF9yjNkHMElQX6FFVQ5PUNlfQl4cRmahjg
649vS1DeXjD8nKXHp0EvWWi6TOx2IZRT4JjjAB05Cp08am1Yeuxqmubq2pbEeMLe
yBMumcUTt86lsjxmHxjEjgeAVZfA7urpDXKkCEKeC8iTrrKQ0GSeyoiYPkT1bqVc
5YvDh4boCC29PnW+6ugDbPd8bk8HhzFLX3HIsWx6zSb6iGl073HHluirLXsT7Ovv
BvC9/Ze5MZS2x5pyRbR064r7f+Dj2zqCHvQrVCt33NUcbF5axj0J3ZUnn+BALD+M
R1OAEM1JNZA3VuDLrI1B5Htd+qdyyjb/2+O5Qsfs25XiW+/1Pw1kk7awY6B4Teag
yinJO2vcsGEWd517PG+krCHMrQQxFnWMpusvDmxzvc35VylBtLVHMqdNg/5BnDn2
tmBmDz9L1it/KD1gtJMfBdQUysLSNJrwldcNq206mXwwxdO2BQZ0qx9ggMBvmxEZ
IjpJGbR0cYHYqFQRBoUvrPt4hLq7fxcAKBjS89xJnucVq9ox/2MdYn+sndCJ42Ii
K33eHL2mnDP8vBN4q3A88eX4boTEZZjqAnoI8Pgj8vuN8UTkD3bHEEe0Jys6WkuO
riEPX3IF7C0g2AiIu5pyxbAre93hljUqnL5igoYc3j2Mwx3n0C7GFgCU89U23qI3
xEEKZxhO3say+aKGt+I4Ro6cwcAUcTkmFw3YPUovxtVLEiFwZ4bwTrMmnHjFquaf
5NGHiOnay/210/+PP2SXVFvJw2luDVecxymlMSXfJICLmqgOYD75KlTkM1icEIRa
qDLevyG0dDm9WGTWr/C7nOLkSsJL1hdzmtI79ixokzIj69nSFcm2g4tBPvSskCe6
gEAFlc+UZ2IfFYA0FU4HbaaCbJVeHDEBMkTMkFQKBq1fqyvhllteY0A5mkoK+c02
wllxSam35tzOThUOxQ8zEu5I+qmaOe3hd6aSHS+oFl3atmj6CGTne874cHcBr4+Z
tFMm6nD5nplutpqy15H59xeia3C0x71MqVpX9pbuU7icN+AMs/rbOTBQ3Edw4juj
57nO9cF/n/pcpqX1Nsrh6Q+qJF6XxoHgI2wwxz6JcRVwcDDsh00Vi4XXms0AD7tR
s56FOwg8Y5mS+BeVJVG2Q5lNGTbX5uLNMomQFaTknkIoUItzJAM9e93mYvXoWQOn
SFBKdgRilRjVlnXCCRguy6IxznVS9o3jWOI7gKEyGTW2mGDe276kVAwq91cEYBAu
OrhBAv+IH12Hyxz4Z0V1TTrwfmzN77xiNenQSsYl1cwIBcCcSV/uIZ2PlJa7PedE
oudXyQT2IK3JsX7i1qpHxUc8xscB+rMBwmlKHO8rMUTY+qTYs17vBd61YgOQeSW2
w8IWPA9WosVu+djDfkLXkdPwpg0ic7FMEhoVKaP5oUwDBt8jz+rdRHng6YJHQyp8
NhdDnwxEcBjcU6aCV88C1tNSbCKIPD1PQmHUMrC/SD8KbWPFV5jvNNb+DaxMxMVO
pZYTfFwbFwIRCqF/8N44AfbMhysdFca++eEsNUoAEOzLcvBXzNTOuDafJXdM3NBj
x6DXce/0g+lxeTpSd6uN75nV9YajyisJMOGsxmbo4acdDuq6hovzEBGqHovm3R2h
11REbpi1IbVf4/2dQcN9SYuV7IFFpvcrVmn333JdPWt/CpOcNl7+pu9r2Y3uOLHa
jTBmJdLOrT7GeEHJwp056L8x2rmzt2ApVcE1jQ+Te/YFFiMLXgyamI/KvwX+NdEl
zgm37d2/IHHWSn/sO0uhOeTlP0wIHWQlw+5NTKLdWe7sSV1o974+psumMFMuWduQ
si5ISeF1tFjWpx/3rVkl0SQxpvPyd4nm5h4ldPmiuZls3/dB1DSN0pI4uodf4/JH
dwPXIu6b79FO//c7VhWSzYA7OBKa/vtaF3ispOomq5gY4GZc0EZnst5RNAi8O04J
V/VTKg30q2li4lG/65nNlxkhEkdHG+L1lAM2a627nXkxBJhwK0g+5T3kyzevRTgQ
tvt/Z2OLUxDNH1NOnyRFLFqGvsR1+sxsBJ3iYnbqHh1XI3Tf50f3iYAcg1P65YX9
Emx6MAP3FS2G7WnEBwDDi9trJhCDueHRdTAEf+/swTXGsEZyPVlLyy+K5yMexy4X
mlpYLL9rh0NUIA09UQFkzIE5vZtSYtXw/1J7sCWqkCJALk94F/XA7TXcQDFrZLkT
V15rXPS0ACftFn6/zXMsVqvTaTPCshPjFoxj04Ke/9qS7TyqNn7UUkLDlGLFedcH
203qGdHcq28Xc0o93GltH0Np3n7OjqtJ8WUSrW0zv7wMKgdgcrEyBfS9uuzSFzdm
Dh2u9EOZcHwKuUx5VxxgHYfORibiyGRkHoc2OrWofKl93qz3w2asgheufTk5jnTu
AY4utf/94waBNkTIno3rAoTuhiY9qZ56MUFZ9wJcQJC4kjrJGHC5NwKR51WIY1iw
xluoYFweixIMaGAOqu+wa6lwgPw0vpCZuMqqw2IT3v/yWhnnc6nO0qB5HZ0OCRVp
xUhUZr44wzrIJl/5kQC1zrCtaHiwRTESmsX5GZBol7I0tb3ygqL6BbVqqHClSFBs
o+2f++/KYZTgQzbVr2sHEmJZTyrHvTRT6zmRJfF/Mtfvw7Of8HzfM1y6kyP4Xv98
M1aC3CysDaaghgrPF4v4bzWv+eQtAVrrGNR9kiG0Z+6ZsI//MXJZp3b7Ks/HF64J
WiAcF8kUi4aypWIAf7Ba/O2hNFJ1fVVtWf8UM+TrU8HKr9kMQeaHBZj9jN4Kb9Ms
TN3mAYkGz8Y4Ps16ceydkh4sNRNG1C2oe98tiIXntwC1OdseTftg7K2Wakp2qAa4
4ZrrsBRH4iEZEIA/APMc+dqvE4sgqVrMR31zRn+eNVF4VRgrqPX+gvm3gv8R0aU6
D7me70ZI0E8s2aAGzOVcI4FQ5i6cfJDKit2OuvJC7lweWDjbXiIs4lMu1D47cpnZ
EGk1bnVdREicJvrTR/kDrjoxMRbKrOyMYKIISoA2MBJpaglVvAD7lOtiMlBCNxK9
zI7Y8HpA6BtSHS7ij+KcMaD3YjU0RgNO/XRqjPWAI+BxVTaZ8KwxaXv+xHLGxl3g
fTn3bt8g7bqENR1ymjonjznJ645aGn/VmeTRFyeBx4e6XyLiPBeTC/xcOfXHEM8y
9Sl1KW8I0xhuTpNrGsKPkKRkhSUu58n3+K7u1p0Pe3zRdXUx+JdqS6bj5zJOPehH
uoXO+UIcyT3DZ114tWVIEWlIhY3gQgmMbLhqLWZDALLBa1gINAY2Wtm4AZ9UqGfs
+bcBUlNqgjylwsIdt8QbjuHIchzjuOjxdy52GV0EyPaPJ/iJsA7Xuv/8FoAGBWrc
trmOR93B6Z9yRdt8hXPmcRd7Cw60Cu0DU5zRwo/toYivXIffNaLgck9ZQaKTQ1Rq
MN3Uv6MOsKiEYma1IapPE9Jl1GZOFg5QfPtuVB0U6xuVPhgV+xebjohhBa6aa/1n
CuCDDOrKRl7q/84LUUHL30zTg/ZckFb5f5l06LTYC9F8f7Qkii612Z3UHu1CIUHn
y8blH3MrozU84em8Kl1r3aCrqaF5Qq7yOd5iQK5X7aPQtsdCUw7TYVNULUzY5ifF
qVKfydYgx8pQhR7fefz04qHAM+J88RBLoJ6WK61uPGUucRZfGvahSeJmsKSlhTZx
K6cKIxw74wZq8IKkP1Yi/WMpjuuyH6sc/dYZCjkERFLvyZ+ZrJhEDjp3SVSBJLv+
5RPCitzCaBi6Ptrhw8dewA9jQk1T1HbrrxEJVxm0OqLZzL9Uv16RRkcZkMdb8B5i
igC3LBNpSqm5eQwFIlqfJkUK4GhgCDYU+6GxwGz2jHqq2M4csSG+AGsLsDpSqWYw
RyS2zr4WmC+nvFeuzUs4x2lqsAB3ug8QuJ8v/B9rHUzwwO9guopkyGX7J1lkelrc
OjWq8Or7ZJ5+cg+ao878FP2I6CEEtW8vRLAyTJPpb21IJg8/KV9F5Quy0t0IktnH
AFDm+HFcoyBP5q03MdmArdfXC594Y2oQPlDppQRRQO7xzZvTpdS8IH9GEhDLMQRm
gdEKiCO0Yyqj5dc/JLNX9mK2PAcW2oKh/X4vuPF6o13S6Jr3Idp4JSdnBKUpuzC5
MLSobpCh7aZwOCeZg4OISmMV3GAefj3BXQcfQ0yYCvGtfF8oVQTGL9IFM6s5ZV5O
pEmk6yXooqI02cyCcZ7R3+PiyTx1d3rHNvPw9KoiIe/i1tNdU7kIHgFaww+RBt7z
TVgVViFpe6ilxwMgwVGwst+ujSfK8TLSLsCWqignPTPMeBML9pqRxBGZqES6BbUG
Oa0+dQCKvYs7IiSXz8dGTiJoj18apS2DrA8e3rOMH7y1EwskaZuxwcvcNV6+Koev
66pXAiM8vpaTEnbnCUylNe7Y8mNqzPA83ym85vkWuJBZV6hPgbJ8nAJKZ2jteJj0
UeLvYfIMSiMBdJbLdpGya2rhfiYwtJJ65oaP5hOmYcBpDE/Bt8Fgr8hYeGRQLPLa
1tDHlP0uje1BVlmcrnBOp9QyXWag+y1q4101WoED2BFpaH5HkfNb/fpxNzllIl9w
QNcec3gRNHPe6Z73ZeIhcTVRWVJGMVaaYAon0hLRyNqOa36eTfb+CRmCObpTH48U
nZsnLlJ+M07MtWOGoI0pxBwOBUNbax0r82eLnAr32Uzy9jOefez6g21ATaMBQwC7
Sr0rw9qnYyCFFjqEGkQ5dHqFA2O6intvyWBjeLLeIRsFFIoAKNQasAm4z6D7nzG7
AKfr5MYIXZ6ic3HhRG726TEop4a6nKeAtjW2Obgb3xCzDEdgjECJ2KFGmoiuS8bo
XIn5mcJHiVlZxTWcoyoPisHcilEwn08ocvN2zUK8jRROaoeCvlSIZ5zDdJKrJIDv
skCJQqJrZDhLz46EvF8tYCKaGeTJLjicz1R50VCh62d3M1wB+J/SXbiMlEJQshQx
c6MBoszv0MW/itCSgu3EczRUSpQEvqc5KbGEnpjGul3eTOcNRaBWHMJQaPPNqQOu
uz2BqiXox8donx3J4CUrPqFli2aHUeFw/AAQOQfwNEBIrO5cdNbBRDBwIRafExOW
kRxLX1waYvmX2zdsdDcB8SZjWBZ8x2nnuOdUy6bu6GYVAKwqpK9BrBh/yyC/FKYd
BtWltoPYt793JdDHuRiiVLWxvoklaaqDAZKD2lseFzyvaBiJHc+Ov4wFAdo3pavI
+FLKoy491XW9x/az1gZSMA2FHF1HD/HT5irYKFJxLL4iFjw33vCfBmPqj9gOAUMC
obo96/ApcUo0heHp4t+e3PSZG2YJc3LctCVvRX7g9fb/JGlKOsfUtKoITyTngRT0
DVXa/mSyN64cny/HjXqeeP/O66jtr9mcscmblATu2kXzFJ9HAU8tHp0KkDMhS6Jd
1LLyqp+3gGy1iSSZCF9ZC1SsBbAxhDFllu9HI6hDDQa6LzPWJf+/3fWEToSAZozU
G5sO5kZa1vLouOU66IAuupJ3p6XYcfGl+PBT335D1zLnRnpU+m/OXKwLnqROPgIb
6sBdjWLLc98ENsOhhWH+wt8ogAm90eQwQypb4Pscilrc8Ff7ncGIGxYAOa4GoYhm
LJZEh9sl1q9DI7GdIy/aDPFMa2Y5+C9/WJN8aWNiOtMwoUAroPQMHL5kZJam53Bm
ihvSXkMmpwsV5X892GTqBT5lm5MEFxTstpnBFs/LWoE26sA/FAQWaZx+oSdfElHx
XjZczS8epvklENiXAcUzw9KgXC7mRGmAhP44NCPrC3kCx0ryDk4nu93zhJ+tdiCd
f5RiVOQUAsDshhqhFw+FNXhxwRt+LwZdxJsMKbtyGWykloIDuYULcGHGXwYOn1U1
fMh7o7GTUW8scc/RyMnwaPLasNlP9LzoUNxoD4KRxKe3szrEFT0R/DuOgcbwqn+a
hBD305b3g31IFbZ56kmnohQ970FaR8DGsz2t67sfeLmsrcOUZ1mvePOqF07Yr1JX
j/l1hVGZHz305D7v8xhAAuUqH1dQFqEBuXfboq/3RDeBlpdghSDDEooAB9wqoDad
TQK7LgJE+9PfNMdvw4QUgLX4Yg4fPIrIyOOdFX9ep2wyhaze4ockszYqU9+vBIM3
SQO3SW8yZj2T+cc6//4uss88PpNrEhjkHf6lHf09dtY/1HwriTZMi90S5rXM2sxO
B+YP2EGOLD4H2UnoMXwupEOCVyQtmSobAJTtuPigmykNO3tyJ/8k7Vcz9Qei7g7u
AlYnYY7hjESAdjFR7J8QCeUAiuOp+aFcMrk62vvIofI3L3U3QnC86231tO9q4Ibf
dn03zh7T43WhyJRKzm7ZrMT1TXjJ3DPILeAOcXevXbhOA4Ll68k5HrdvFqpV+VCB
Smx8J9ckCFYmvaCtXIAPcH1F8my60DCw/ElOeBq8YYavGTSHjcOjGebfh93StHlx
T0sVPDQJjS8CK1WF8m/anZ7jBRVHD7NJ7kw4f2Ond1fUJbzRg1Hpkkz+1yGSxzX/
b61wYDZigHqavP+hN0aS8A==
`pragma protect end_protected
