// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:54 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
TVEK1QpSavgeXOjQYwb+RCpCG7aSF99ub9SCsHAYyAAP/lNSp+Lom9h8M00qfs7A
RcG121AXPXUtTkyjY61GOgWB5kJ4cX06ElHr6tdeVtsw/78kwmj0VVSJFcEkntmy
qFmoCJPHuLldwNb2Th5inup1w18ZoBD/GKTCJLr64/I=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 16992)
RX5hJE01k3fo3CAUT/xbebtdnfbNs+n/r2NdDqytc2hgBbdWq36K9yEVc3os4dTR
nLjsGaXzf4hNuGQ6N8XnXJoAbhvu9QVp0Nloq6YG8VjxYdbru0DuH4gndTO40Ja+
NkjLGuGqe9mLGjBqMQ4i9sIaFv/A1W2d2xPjXUbW7ZrC7Sz7aeY07LJieMWy4l4v
hg35ydzD7n+UYyaCRnqFhw7rkyMHvfHKTSbX0Tei0ratSGphcEtdXwsMMA6CLV6v
IyJOd6CeKtPoTthj/yMVbjMXqsUno7jME1iV+sLchQqazNDTfPDxPYR45XxJ0iLW
BA/Kb2llXm6C6RuCCxYhOwu/SsuTolSP26kLeCi8MU/GJsTWXCy6IUvaHSHSPcoF
ZVc2cK6RECq2D1xfRsIzz3N/pi6N/SXrkrVIFGC4O+i6XyXFAMyMb0oIPXRcy6YK
HARnSOReQkM7lPBi5hPGQipcac1q78FgzmO6D3gLF7D4BMfzlEc5+ATc8QhHWRcX
eSRUyPO7TMpaY/M9FYXSJNrNHzkng1OVulpg4LyI+Co3CoEQpHRTB1bMEBHP5+Zb
54exHsyOtuPUij/gWQKaQhHncv13tH5V1kEgw8DQF5PfwKZLmKHIv4+4TsLw23cq
TRMsd53kzc02Uo7gbWKb2soC4QG3JB1izLOaQoQfObc7m6AXKBY4EtdMOqkDhyE+
b/YtvLVFrfv3U6hpo73ZLC1i42zHzr0riGvSwcekKOoxZdMmXPyGlIebIvN5TktV
kWwAhBiJNO88jab3nYbl8J+EzP9fNhfH1sygJpLE3PgMmBYUQ1j1RL02GfLO4zlU
3s7XU+lw3NEXEoi1n0wEqLoUCSmHSKWQooqIWnH0d8pSbJN/20F9Oq9TGD9Ph5dL
Q2fMejBkldbNQV60i/WumNS2skWmb/a4uQiF2bzTgGKrX8JUw/tYbiRGMeHCanXV
lPSi1Bq3k6Lo7Ph9KHhY77w/4wVeH/LJVP/k6AvyOcRWenB/yEGMsre6HcTUwwk4
UM0JdBNwUV3tkXG8LpO3BZXOoJjeiaieEJhoEhWM3R1AMqR2v3JsYcAWdkIZYDr/
ybcRGMy3Sby6xeKrIcsZ3FJwIc8+pgLu9EeWT4dILGpqQQzxSOhTK87I3ggow2kH
p0JTBW8g1ArEvO3yIDX//6X2ImVTJC5mCnTtq6PMYotMFd3ZeAZih7n20LUyh5ZC
i4YzBWGLpfLASfSPRbUJjMCymylPKDfnLxI+VmbiO+hU3jy0c33xutTk6ynv5/IF
EiXw0xwz8e1DUZb9Ck6ZJcJYRHreTvuExyMdPDyFmNtSE6J/H/As9PKN4zil+sTy
QOQs49CAba4SIlRPhQp78MDXLe+P/XEDiL8kQW2A7tn7sH7ymSrBErRRfLBuIp6Q
2igtMO8M/ibtvl9jd9Nrk41oXfgjHQ7mzmmvmJ43xZwgz6nHsUdqnz9JfQqlfrii
FrO4RvtP80n91hGedMw6AQGSaDkrW3mHG2F7PMgS1boMvjcriJGbdqWyxvVCnHQZ
WSZkBYm2KfM0jC64s6r9PKzSgCW4n23cRzNPJ9HNtPy+aaqT6AO3b6vWAq7LUX+q
4MUMczQPXPF+VxwsDd5kDjr8NXz59DxHSlCl31rKEjuT9+20Pt/ETp3be+nRD+RN
lRww8bHmDtdMz7uLyALIIvCnX0WXwQZ1Hut+c0IG9oxmTSfAN3s5hvjePYCMgsNG
NZxJCUA2xMd7mT6N6YpWQCmNyFBXN/Cq1630kVX5hr4GZwyGXZ0kUq+MxPBfLU1f
xytVR2ukwd4bfLSvlatCeQg6X1fy8xNvtXuG4iTkS1Yo+Ng5i+DJjVuwsFQhwXlB
y+xhfMmOhP2bzYDRcDdb0IdE6m2q+DFdRbdE1UkBfpzIArJmUJ9LTUC7u7MljYqb
y76exb1q0mPlA61xMcfSDCyAy64EkobJSnun5nwikY4SZpo6HYahLy7hVaSIuZZn
AIsJYnJY1IwLG++KcMF62KIeRa3URZclZWBR8cQ/zyRrMFR3Xffg5BJv7QIRJoHl
nDNGbH5xhO8Ah3eGYakRhZD4TM+mNk7XZ8K3kBbcHKiWyob+8DXTU58wzv98WTul
ffuW86l0kslFTfVMzVwuWxoOAy2zenAu3c6EttDpaeOvMAVEuVWTvMPQol2G9Tfd
j1jKqlwXHBRjoExtfUnWoyF8kdtRdenTmYH/bJPWPeD6nSa9UYom8F81INFV7PNc
pT/GjjYXf6PHWVQf2nAjyEyklAewbaU8xl3V8C/yazOF+UAXEJqTBMAJc04ypkgN
p/mR2tP7a089jOCPNxhvcwgbLhXp5VtI9mWcusRR9WiEgk+wtBfBV8HjbXIFg7fn
ZxyP/7ixdaJb9DXwebeYaMnslHujn5nbUXEppCA32rpHQBtkVy4R0599IsuGChDT
DF4nFKo5c1+G08tCqxISh/PRo8QQ5Af8LsvwZxO1PBYben6ufsFtBdFMPC5m60LG
T1r1t8oYO1dDxCz9JGhenFrsRIQBPO5Sdex323LWysxFjzNU51vjKN5AVFJ/Qt73
LxuB+MpR5iChklCq8sxG5BpaeaOrP4J8Y6EhAFRxKhmx9uHUpUU/Pd2JFoWar77A
K9r7B9GXQy59SjzG8pclYuPr+EPNibQFGMYRGXqJTJUOv7gnUjk3+pJ62t5wtZCL
rbxHvFoz8LvaykTSuQPtLGBzH34kQQElQD2m0MqRUG/7lfqPbH7aqhCaJp2Z/N0S
5w717Y4YVEUJxlgxOCUM8d6JB0MwwGAxzCZsQuciITpJeVRVyzpTdxI8NCM1D/ui
6aD/IrMnYOy/X0L3qCgXq+cx6wm5BWIE+q7E1xr1IKhe6QaPHNC1QzyaDNPlfcgs
38rkvlaqInG0rcfaXLDMN816qImoQg6bAkubnsAcCNLZ9uHlM7sqyeTw/btbYRXG
UaI4XwGCks7J+tGopclT0ygWyGDTUojmQLbk/Is+MgAlVrTyPyWd2fuovFS0nQio
/dukVJvy/la3DC4yidk5pGZ30K1rYJa3ID3ZDnbM+sBivT3ZjUmH2NqkVAYyaQzw
imoWLZ0SG2TxpJJLu1rXzB6XBMAuSGqCNIVTKFZJMUXquspotYh+06q5ie2zkrLG
ESEZmdp2QKCYX2eMoW5DqeRvRYEWZ4vvysJ5jHyQP9dIoNxdFIj6l4WaHHiGH9BV
18zNPirm/Mwuom4eP7+NnolMb5SeG3zX5+NGcFGKz+qmr7aBZte6fZVC9U9a8gfP
W7Knipp4ztSFpe1QrUtm7F88Hsq8F2JScvATFaI5CXjA38qmz0xAkJtPmK1pxmXZ
oswfbH6GRcx7kAgX2Z/6VhzUzPdDN+Bew5Z+pcvX+j6Iw8tTgv6HkyOaTA0bHdze
zptLP9mCWJ3BW6NBfc55j1RgVCSslX8V6NO+SIhp9MEipS2e/qLwwQ0SVSyeSdNX
3pdWkP387nY1N1nQ0FUn5LmRg/OP1hNWmaNg1WCi9RQt4e0yG4qYNtZqqFbcW5Ow
Oo2gLJVBNRLNzTN5FYxsCthk1tw/dHblVvJaCmOdfM0H4cMxlD/eZ04zHD3tOE8V
P9mTn8BCpZXEwNrFXvSmBU71VXBnPH3rGzr1IphtVQFLgt4kHMKNjARHcKq0O4xn
enFMXH9Uk0SmUdptES4VMkwdz7IIl6dFMT4PKpeUixhr1Fyl2fkKgG18FXycLwKK
WAhIBfQMVoxbNwL4nMIIuIrbzwESVjgNsA9h8FmiRkqw9XJx+DV9JhA5cOzuQx91
LcNhsOUIXPudk4cs2QjEDevrX2Ot0iRzZ3fMMd/H7PmDWlNJiq7vwLR3HRvS2fY/
su0rOZ7LSbUCpk52odzNLP4yp0Si4wtsWdysScKvv99gYUaAi3w5j3gKsNQyWOxK
p72fq7b0roLWhupzG/PDRTkxcQHrkn99e3pyVq/09moE+/44ZrNKcmmtlfHBvsrS
ZnzrOaoVEV2hDLYy9VNzEa0EJlwzaI/Z6CtIPxgAFHTTaj0ANrDLcerVNDGttq7p
3d6xsny+DoxoFr6DobyBcZRk+hCWAR9PJXRUgi+BrM0LIjO2PFPwlGCxBPx3h7ZM
Bkq8GGrBWvgkwC/QWdbafHMdxgBDfpRUu9NUu4JdttX90NpbzNShtAkAp9FMQ1i9
//9ourZ4hRY1p55RGSLfFsutrSdbnPi9IGVfdHrGMDNzcT7zAcBuOE1v0dEy60Jd
kW9nhDb/Fq8uV7XbaaBOZYq6gqN9w46ACbnBYCdwgYtYdq7zl9RH5faC/Us8HmIx
ZY4ZUbYqDUPLI5n0AchRaYjs4I9AWH7tgt3Ie12DOU/3HtVYb/7FALNULFjh0u2c
hhU8NflzmBx7HibqJmmuvAc03UQng/1ziFFaXGPqRRs5BwfLyAmLvPgd68kE3SFK
zxbgL513LdReu2Fz87WpLlUs6NXeaCKtjeRVXQ0F+1S6M9Hwx39vSjTMeAWgQhbD
12agkWvlkzkJapubGAplNaYte0pxrwaxSDqTymcMpjbD+BYhfSIQdV6xj1BuP25t
+Ar7vRl2h1xAI4PSWIGf4S5ADNTKKGgoB1tIs7oi0oxO4JSJ6qlf/73H7RI3haMK
6L1u1JQKfGE2TNx3eBrkl7Tx1fRJ/KCqzCWSc9ttxf4fDMhBbhCwCKyaH6V1qLiP
JZ5904Mijy7CjYKUjCQnAxH0qVZ385GZEZcqQaozwGfxu8Z21fCEiAZOhbedth3o
KLCougf2SotIQJEOSkvM7ApO6hdgo29avXL6tVPhWzsoEVvk4TvvgajOkQeQjL8M
MHmJFKHEoGACeP/bocDKy99helwXWcQQlnyF6sHbDlxxyVnMWoImJx5D+QdEiX9g
1PPARfM83b3PhcjJx4OhsDld2F3iwjJmXcjm53sjy1Zws1tHmQBWhIARusODYm8i
tZovDL4VxnJNi2VMHQtuIzJZQ4+yOleQfhPGIX/Xmq+ea8cT0GmQWpDQjhfSVaUI
dOqsofor3eN+L13yJTqgiRQqMAyr6FD/zdXYiOYKX88jWNNNC3I50DZZrlhq15y9
b3xnsxGONm7NEEeUZl9BW9HJTjXIZICLstSBG4l0CH9x3DLvCeP7jXo4PFaUmg0F
5Z6NKFULc4e+Xuf8qWHiP1HGfGZsu4aLkmVjPHmWOUaPDBMwLsOYSFCj4JlOFoX/
TGo8z997s9Le5t1AFdYwQtPkC3PwneBAqPCx8gu+84nQBKH4piP4mg0L1a8brVyG
UUXJ3vXOM9ym2Ei90FE1QKV+YInmCbViqPZscqMpElsxFf/FsSvXhpgHgxajoD8G
hXzaMDL66KmeLpwakQlv2uIoAO1hopp2+62t7R8/0n9jjPoY+iY+ZQl6fLUipPPo
cJX1aSdnryjla505KxoDVT/Pl+sMp1X+++GProyH7Nn5PmCvP1T1Rg88AGP57NSG
a4Cc6BaUQkVNEjeo5qjw4f2qFaGQ0JpwGSGmdqYsYuEtEDH9l0NS3L6exCr6/536
bchquZTkYXe20gqgMdTLeD5r8HdKL5tx4r/ETxzV1tNknwN4nFGl0V3vxmCVr0YW
Pu91JXwJ1T4De8LTGYtrkdczJ1aBTn/rby+fy+bVbtBukcnIExPZBtAqN6TfHjTh
Gh9V47MVgADkDmASpfg4vDNqH1658UDROMxFZEnzuCs3SR9FOOeV5/y6OH2Qj2FU
wSL/nHRfPuHm+M/4+cCV3lsfo8DFv7oQ50uWIz2CUGSoxJDp2UwDIsZeDfvAIA2g
Oio6B7OdPvy5AHCvfslmCN/i9km8yYvR51n2syJlbMT3tZqREIeNdP0yrmGh8bAW
0RC3eBajT/gFRDb6HZ9uG5q8EkDq5xYcguRE/gelAkTaV/4zq+b25rLVeJy3Oh8d
hatKoffwwzBFsyrSLLybYX3oAM1G1vUByAq8qH3CaOEeQepABH10ILLqHzTw/nLd
yZDu4ZcZAd3sgdD54YgRHZHVy3y+PBfyH1o3py/WrGp92jKj5bpgit0bLjo9QGD0
s61vGs3E9Dr5LVTbzs2jAIKCnAH4NleEZxs3vB0BKMp6dq6ZloyDi0+OwB5WmdkR
8v43SvWdYlZOYy2L1NA9xTvV432pdMdRaquuHOl5z6Kb6baGO3wN5LWViuxBD227
Urvmh7Qy5OoF1QVI8qHS1PMYODgXGIGzcAl6j2kjuOoD2niYTwgi94l5qkPYTLCX
EKAV3aRy0Ix8cxMC9Uw93MWwGmEINcJ43hbJIu6r4IXgKdxX1jTfzACWloOEdMja
m/Vf6+AMaeN+byX5l48Me3q0gkLvGNQWk8biKKSv6nhlMiYRzk7qjvvLvDE2l8Wc
9Ke7A2z7cTJbOBaV4kbMAuGdDKfdul3pK0/Yvag/JPYrxYCPcjmYFWpxWOKL5IKU
jQecxDBv/yzu7Wto2YlKvafiQG4xaWYWl81nsspV2lqZcQCbO1qM7gQ+5XL7Y1Fg
0y2m21c85dsoNqsr59TMq9xhdnACOJlZDwfTprN8rRSH3eDpwECQ1F+EIntvPcSP
hBFNbcX9X4SpbsKp27aAl1BC/bq3Cefd7Q8RdYnfowzES2w2kgWqXLtj9eYXEVY/
JE33nagl4arQZNnJGqR6Iyp0ye+h5aKW3xyU3oIyTd737JCY57B+JOs1A9uhTsd1
nCLYcOvYTs+SsPbCcTMDiXFDhg+qYWZUIRTJi11W7HyZhoqmzmJXD95Vq1reQ64t
EOQ9FPIuQi4h71q4wAKGjZX2BSAqb2bqyykTuyKsh6f1N4WZcrkRTLRyTJnKt6vg
n7b/YjZT1TdvYxE44BtiJNEKiwI7X454yt2uH83fVEKovmupTCxVQrPcy+oWJ14Y
6kUMU/GNBOH8ALQaQo7Mnoz1YTiU1hd+1czMzX0/6cvsuoXsgA6RT/GGFQRCLLOo
LlGgYdFbe04O+1jmHRA7Hvu0MoBAfJqqs5i63ujdqD3XTRqoQSzHDFV7eQ8U1lJH
4btmswZmhuRKjFX+H2dxx2HImCnQMc6b2bB64t6+S85sWTR4ciP+341NEMyRT/gH
f8ExFk4wbxCs+TCkVnFl8WylB+eQN055BGLHc8o8MJFYrfXhfyhzb456PW+1vH6V
lkqlhZ94Xwaprz2GLhQWseBs+tcyiBC9UKEXAX0oY9qiG4mPv0AwWaH/6pMTkq7U
wilNS0Lllaw3VjL4tys5DU3G9BS6QweTk93VZlsOWcLE4yjCXyy2lunPZH+X8gxW
2oXjuBryH51s9cQw2z3UH3R+tsfWGi4/s7rst/Xyktmlx3czmwwprK1/0+hiHHQA
jzSiGCgsNB4PE66b4W1r3oME7HNO95S64jBRScAycsSj7fcl+68neeRQF1Ygj405
f8AVqaDAt5Z9mTE2buIEkasB9EGOBgMqhA55W8S2W+DH6ubgyEqxEBe5y6G8sZzf
qMbKcSc181AfzPhcueC8qo27gyCa6XSI4YuJWwCWIAWe2EgQknDNWbvG/mVlbdsQ
w6vpGvCf69PxacOh2FzvXViWjCB32TSfTAjShPkacTQzmXf0tnL4SVG/6vjjPnmD
9HH/ukVZB/6i/wvmg2HpQ0tfawahOS95BKCdD2dKED3V5MR3NN3APOrJsFQjkFhl
TCMSKUzyQslcW8DGYSrE7vzYAo9QQA6yXyAx0Xo2qLII+/72JaAZ+zfGpYwwkqVn
D+tW8wFYSX5FhoDt4G8lg7hK3hnFV663K52Ji8p7NQx1YMlAiufPGiTV58EZ/GzM
3SSundxptpnKitp+2FtCMRAN0UbYDuvKK1n936HRXSeiSYnfS1I1PIv+bejDrjK/
9om2e8nG6TtLY3ekdetYIfvNO5VfvGJcyB21GvJwYp2sGZSihAfw9xe0DtEdjNav
RQEgWJ6uJ46DhZOfmttuUR+cQQwqLpmuvm8NZE4aTkredW7ORNFggFzn40I5jS+C
zbajSAYvD8DISCKbgbqixX1AFfhFocYweVI/WllkhAKuENO4ZApyv8FEt1EN2OF+
Qyz7R1KpXy9LhlHzTWHLwOwJZiai9xRkOOof06pXPVIUAi8UDa3wUX7vDJlrCRCV
fRu2zyIrIlSh3krck328D7vV2TbVDQu2Zia84QQ/jXeJSfOKEZL8YNZfkkR/NasQ
9OMkQHex6LFIar4kD1pZd8b9AYSnuN6Pd6gS/RxRbKdfMbZea2NVaUJTaE2D2kN2
pqVekdC87ejM9kQ357dYC5HSaqZL+wdAvbutkQSJ/+FmUGGzJxCbHe+p8yuRj+c0
st/QeBrOacCRrCLM9OdFWQEl8+bxAbOx7NTBRwq+pKRoNyxAw26wFPQUmPBdvIxt
CkDa+UKvGGqvguU944BHwazxJzNYlLmA+9phZ6esHr0xA96kWaZpKbKlzFaOl1oY
WYAXO5l1LxI13/c8C/Pi6e7mKi0bj9IzOjvTV1LMyda+dlRhm61wEXlKoX2BWvy0
d36MZRmyWr8L41+FlOIQY3b2/JBmjRbFCBFUqK+ThUc7dmhBrCI8HZ6sa0pX8FF4
+gx39dVGvrdL3ftl+fqCoBZNSmR+tIXjmrpF37IBJP0CdLT8eeGlzcaYnS+Tb+yV
qloGK8I9stivZqEaSmSw1c5H0sKoFzswWM+P983r0MC2TEMp4cnXxHN3GFLYqX8T
9N9GeBsQ//38DYKIAEzUNed1CTnd8xUr2UU7/cPxbD2SrUs4ZqW4KGy1cFFM7dyg
0ZcT5piLuJl/9/b33b2fKGFQ2JnDQPj/oGESD7EWqr0SuuYrUj4aj+XYr8Lb/9M3
mqtGbGvUa1LlCn4ogEmmj+UOhl0Lv+CMd7Fq8T87fiKHlutzoWcovoF+0d1DUG8u
UQiUY4xMpd8x70iCnSPMscMPhx4y2r4f1IxzMoM7Lnqk6FaE8bZjjt9xBODVET97
CPSiTeJCOx8+vvgXo3gCQ1fzOqrel5Y7BI5m7yOdsHORjaaH1uEzy3hMm5Cx5pI+
tHT1JripFQDewvbkhTyz4sb0iM4rtH5/NyZWQTCyFgrsayRMNr4FxjWAsBVFROUC
R9Q77uyep7D+bZqpPXRkkHsjUD5c39kePV/Uim8OADZC7EtXIjUHg9iO1YFBm2OI
khP9ML5Aae8t2a5O5ETjcCIWcUZdSBe2j3WMEy1a0uGs8FTnxoJf+ZWRoi+VlG8L
hLrj931o08V5L2yjK2mQajG55i/WnqFJY1ZmSc9afMTzNwaZ+eAQJRtORuqqOEQ7
+bkp/WtJUryPwA7cO6XvxltUVNQ4F0VHkCd2nVXpBAH8sQ3QO+kc5ndocBOcOSj5
EAGv9BlWnJbRzd5pEhX5GclqsBzLBQW5ITP6Pwg/JX12BMLAUGhQwTv2tlhP5gr9
2HpJDNv7VEX6NwlEEy4xOBJXgzStzGv54ZwjKT1wlPSVaxhEXWFoFC9JVbYlQU77
H4wuWucgH0G+rB3Im379diWt/Yl04rTMi1cX8smIBp44qwGqqyPg3FTqJSPQrGmz
i9W36NbxD57E5u/Or5g5phjVCtHN8klG6o8I2jdZyjqwu+w+1a3lg96TWb1FZzEc
hzjZV4G8QmreLNAAGCCsT/NVpFeohoSrgOaStq6SpUWW3FWjw8RMii5npOkxX7+A
xJ/INx6bLBFwPKMj7nOjvo34hwMIQPsXVhrlk6/vsu5ChmHKbHgO8fQVPZ3nmspg
VXUAGUqOpqtbULoUZo1mrbfSTdKkG6uCxgdPww7w2nUXa/o0Ct6gVv9ytNvLmrpl
xwnWw7PSfISeWda99snPkW+W8omuLTXdEyZ0xwvx0ASsDMg0WkOpeKvIdsOpvtw+
zK6zq/dhScmOylxIJlVOQYlXIuMF8ph90KWIM76Trp3jD3Z25H14x9WRfCkLcLur
RIoO3F3KwakdiND5SB7z8yTD0D54oZWKKW8ETMAFCh0Il4qkm0ipadJtHhzQc5Tr
osJyxivuK4OYPwGgCUNc2ZVRmBgCqsuN2ZnrPwT3nrO1MCgy6ofshb1qV5QyMJ8t
G4CGUpIal/Ibxrm6aXgdqGDwUDkt11pcweSymSi5HaFEe/YjTX/JLIj9AoTCdOpj
6Wsg6aNl/eWaghN3UXH2S5J6rn4may9TIBTZgkJ9HLwDsyRG7Fhs3QWtqsx+4jVb
huwig6eKA4ItC4vGn5Ysm3pHWpOYo/6AghP8J7O4A1jcTuw6e/Eu+bhetglmAxRA
KI3zeyUwlMZywXv3amLqztF0dqWs9rcNZr1rGtNhgVQl2VbShAVp7XqLuTc9a0Iu
kzlTC04pknwOh3WyJk+pzQC941SMIyXFzZ6PEXZvLxWW3GR5CqdkW5bzmQOYVubf
xs+ljAUYCFbjHyrPK2vJY2T0+NZeowddBmUUJWlCG+R+bndaGg0Y3Yd/auyKrbSJ
m7gNdlswWM9JSx7rtwRdfHLdUcsqiLaaeedaGfD7kxBGQNF+mw82Cv0eExO25a1y
QPb0HxmwZjRwSJHuxQBq9qczZJ807FYG00byfQ9fE/Th0cTuYAQfOzlGjf0J/aUE
Y5VoHaCJjBzgKz90At0IW87VPLaLhv8DMFVw2R35k+gnolxkT7FzorTwOU/mtErL
cOF6AeqfpAGSFGdyXsYLmDW2R8RE6j7/BKQgCWdqqZRVgjjIJq5Momfe0xro2JLx
D/ZauJoT7ZoCM/rrHibtDBvjjavZUWI1aHwiZ7uKPDMaNPZN4mpAagg7TsCpFQsC
+lBkvPnVhZivjbysJHx/9BQ5Af2Ke7w6x8dWb1RaXrHuVvD/kUkDJ6MRnf+0TNQ6
keJ/BI8GFWAyVDJTEqwwnUTnuOFjl89i9buxpNBNXJyy5IHKwf8CoSSxwe9IO0hF
hccXFqNUHUJ4qYdmlg0YnlnDnNsAuOwwB2t31G0n7tkOlW7ttTy7OG36WcDqlIKM
2bFEPHnMOJcTvdo/SeJf6i2mEuI+NdeAwHBROVmCqQcC8t4rlHhh1i68dypCKyih
uniGU8tpA1z/FpIcQCDVcpsaJQlWPwzvV9xqzw3y4zqs+wFdFE/mGoBrM0iiPSrY
1+iOBP4rR2ACUHlUY7yheCy+C64cRIsMjbuXA7W1OeNavSTp2qTdPdpeoZdoPfL4
OSY2Q9VhiNQy8xysB0aQMhfwIsxcBz7Ia5dtCJouzhkf3LnfV34wL6AMBMI/ozzR
WMI/R63nTxrKjlHJGdTgoR9yAAxX+/XzebwuwjJm6FDDsQIEooW1vQ9VL6/eUfbt
tDgCsQe2YYEpGpmO9ciAtlRXJ6Sh/gKMcLz/rU8tVeX09YDsbY51Kitu3WBeEOkA
7pO6G4wqe4C9gNMBbazGKfJPD0bUn9XrILlivsJU/rHDvPhTSjKuikNt6fM2M+8k
NxE2H/RXnCxqG702SVJFwh9RS/VbSsYFzRwk+BTZZn9sJMKQH4OCMeqaL2I38rYd
NyOn9eKi4Eh3RPy3Gy1O6YoSrlr96qyoN+ND1pCs+wwETrNFiTrUNeqJ0ghr7ZWd
TiJNlosYOVPEeNRnyJ8sgya+/u54hUUCUWUhqm7wAcXbxIIH1e3JzPY/MfNQssyG
bxinFNhFHBfSAa4xEYRZqNWehf6G0enplAWDY2MXpx6cpgripBXD4LoJkylbIBHx
vozbUblf9qEmEKvjTck8i/yFyGCRP2iKg9Xbj/eCwm8kkdJtpJo2p4PSk3fCVo+c
on3DiAi7+tDS3meNwC5ien7Ju31pxMwJmJm3K+X1qlngZwRjzzekVbAclwvZO0jy
Fkp5Gy65K84PYS80W/PNiADd4KZsglRRULJOkAOzFKB7m1YaniDWL71GlSuKWi3a
D92+oTYejj1Ip7akUxSM41vdXqVWAil/Gn++SGaDXn9MgIw0rchWsstqCOrlOtUE
/fZvVcgAKQ+u+pmcxOcJiO7t2E0oY52X3WRXa/JQJ/VTTmEOZqfs8mct1GgMBS2e
L9E3pejzj27zcLsfohKd4vtADs9oRlMRDv+ofMj+X2rZPJvQM4mm2DFRH79DU6Ah
r5Gc9i+nuYPWTMcGeqC0HDbzOA7GpKt9hV1Q4Ru5mBGbNrNaSi1CRBK5iKNtqAtW
K7GmHo/qi8BNsEpGB2mCeX7v/WZ8QC7Y1sC3VZ5qXUf5jXCRtAzEbHOsrAW6MCxf
RLeILF/iYSq+6m4JJz0PPsZNycieGjPAdDJx2yWpiRDaakGgjFOgnw0rZ8sr2tbW
8pYcYLaVXpHyYFxjjJNRePaxuopNIM9PbZVN+jhmDlng+kTkfpPgfIqEx1AWuFr8
KerviGyNYz/BwP5rcy3ITU1zXdidYoPHoMMJZl8TMGz0OxQ4L5N58koMlUqkl5vS
0OCdoqxcZ6ZZy0HJVc+woLKgF3RPqbIb1jmTE6d6Q3XUem8Rk0FR6Vnl+0pgk9ba
kqdbD08pohKlwBC7WX/PdByx1mPaU151zAVyF0BBStbdJKDy+SEpWfaCkgDxBEV6
dNPgh+Ta7GhWbfiksGdFW9AsYtvQuMAK78qUL6bu8mb/Opy1JAIQrdwu0ZxEpEDF
JrjXZ1Vtl19W/9/cv8tU2OpO3uwjfyBLdDMdLC8Ln2LxtkK4hwEJG4XnWfD2fHmI
VxiGcW/DLy/WmuPyviTOmNKv/QtHm3xMHm+TGCTn6SWbDHrxrHh3rSI/3a1z3E6I
bTpkwhvfYPkOYIFNgD0gYsPQTn+eZ+ZYFKgpxmEaWuUXNERgOfzwLCOii6e+dKu8
B9ZFLSFgFCPv43Djui5LgzeFve3ROEBTsYyraEKrTp61REZS7xcPulbU/vnQDMvc
I8G6MpdJlztWVq6Nwi7KWQqQv7Dio4y+SE9nWX16OwKecNeFMaDqQ6ibSfNr1Hfg
8LtpSJezxEZidETNwQocjyFr3KskI8Eg7eCcY5xa9mc5rVGF/hFFCUd2eZTowoCl
78So1GWb31G+0vx/qQfgQz/uM+34I2wLB+WMFnySYoo67rjRgbqxyAgGTWRtJLrh
De1n2pZTYxe+h7ioLtVoNwFsZRRGQFb30cJLP8flnTIU9aUgk5r1fDelA53H01FA
lTaQyAvqAf2HGI4gsyE9qtWx6FG5lJFYo9prdCm+Ltp85RUBVXpMID/tVNWevz6v
u2hYpwTfdDVqd6zNNwwWxpqATyGA4rMyBrB4WniMBKXP894DrzG2yGi5cNQUVOkh
46gGdzneLa5oLLQmrpX1Yt03A+DUtiWqzRYlIDuxSMYtHGBOJQ6z2Fc1Dmej647D
UBTmdmV8niplIGud82tzcLpbbccLMiHwZ++nIp9qAUmxVIrJRYOTyz+lzq8iaDui
nrwZ6XS8SIlyL0mCTkxSF2JMwm9wNY5v/wx8hqBQdaEyaR2z+39MsOLqzcWQKvYM
rrXVSTB8qTUmNr3bPJ5T6hcSFIeqwYSUPUzEkBtGw7wDOp2b6cCQp+iMCxjufaK3
u2ZcR6g9/6iSnK6n67ZxU0TxXpE2VmmF9xDt0HLJWx8Xmbh7YA1Hrc6nJZ+XF3vp
wizRhZAFMz2pB8xhgzsnNzqDcHI0INCNV19H2CXjW+5GJy88FrXG8X6QDKtN9vKq
2LmEOeqfPSWru/G4ELfgdkAEPnuDcXDBIPOYvXH9hF02eioDfgVWXTna6DIV5hH9
+HYUjl8wab6XqkYubg09nxhZzuIC0nFIcUtn964AA57pDjWudxf1K213LtpzzWbN
cPc57I4kEIGyPUd2/Dbh49nr7gU1Ysn3cBek80jDRmUQg3CjvleS7s3UhVCDseZv
YsaJMqaOKqSMLivy3YYitxhGSUrVni5aj14Yf1XRFqyr0J8oU8QMOvvpHWCe9EJP
7Di03417uKLZZwwHUD6eYj/t8e5EvBd7K+9pH+uGOJbRhKPxDD9XdP5MHnVIvfRV
mMqnsMA3/j/CLdg0RH9h7u7DOwGJAoIQhqBmXBKaCoJ1nKR/NRt8F2aCZ4TVO2gd
WlcfXur4l0YISZdglx4SlhrGISfMrZJ+4W8k1NQbhZbu21tENfHnoCii2rhU8BzR
urR0xiAZExKNTiMnH9xR6WWTp5a72I863/QTYFEDEmggORBrUQcMv3LNZ4lfQU6j
kzTnLJT0mAXfZv7ffS5BH88T1vV/JWr7WRpb2eoQkE7m0rKNozuHF85/AKE3UqZH
Cimhfu6AU+3zLFrWIdhXAarAwTIQpoYZOkxDItsjrhlt4omvQpQcQPpSB2Euh8+H
wWu5tmxwTgX/2oqJF4fblgNyZLdKwTBBQWKj41xA2SCqkXsqxfdidRd5dUU08AFk
qXjz6a2v/w3ytCc5YHtALM+iZ/4GWBw4ufKopvNTLcJUzitx/sZKBr38oEFeP0sZ
2gXNTZ8Xsn/UfDPjP0kBY75161gNES6J8lhzT/CSeLW2YEXHPi/nwHmCvG6GCFTO
M3PSJ1InnaITL53bJuqVtOCFzBBGHbZFUEjN4JEU3pElOYHk8G88K0MbRnO9AfZS
pmuJDJo1hCttDGaJ+0ysyKHV9eAOELy0Dh/xDI3I1/C6rhCQ9+UyydTUKY1O6MCg
uT9bDPHGGAofa78XKM3AtQ5UNKqyPZC2YAshHmwAGZOFFgjfC89QLUs71WAMfSPl
0Zpd/RzrFWvomcMHbAFCK1vHL92EgBQlmf9juvV80JRmDq0Wzhs5+LEPsq8JzuWD
SB/ZXNnR6zWe/VkMm0oDjbeqOa566z+E4HB33jnPv7QP5W1xQoZsqqsaqYXU4Bqx
crYKRz3aS3LbtW47Z3GGxbdRhqsdxpXlcFW0/hxWbDNvyT++AnD/J2jLgnO5Ziqa
jCdkvnJMkHlq/F52Qidlo9kVT9jWUSAdBbSeBl6+Y3kfKydbt6d/k1ZMXzCOKE2+
YWT2aArfL9Sm7ROu8H6CrTYi4FQP9vqi7gZg/Kmee9YopEArEM6u4lGBjL764HRG
EkEV/orhIe0goSpddqHwdeXclJOze/TzM82OnU1alk4aQAGvNRK7fJrdE6E+tND1
K15moXcu+ty4VVGhRBh4/21/lF0sceTPfAJrajVzIkQbwnC/2SQQ3aG0i/ibbz/r
lWf8hiftzFM370JU0aZo+W5aOdHW9Gj2cFoPNk/++G5OEhdD6TMm0lQ2uzwB0cWs
QS+g/lNfEK55U9612fbtYKbzHRcY37VY6SKaMQWjluQtvA6ERh3QbqmFXDiERvvV
W0WUiBZkHB12Ovmqyy8xVedHsUT2xfknjMDYk/65WJ5mrpv07DAi5jTLuy6Yaowe
rkPUSo6lHth/79hGg4FDPJ9tRWZiQhmT0mMlS2n8ggqcNVOsAnyZ1wDkn2aOfCRd
lvuj2bZLb3uoFH2lrOypuqlECv8Y7QTTnh8vU0kR1x3dwesLgrHjb6yY8alAPT/r
kQnZfyRyu4mi2o8IWV3URi6wP5QawKNnzSNc9Guvqiu2UjauIoth1GAaJ5EB06Fz
2niiocv982GNN/GLmLVgVPTZfUGELbVIYBWB4+jThznyM+ytNJ6oSW2/mcj6uoq0
SDNoZPEmQHjlEJWdP3DNNR1OENmMKQsmKzBlRcyDpgk67T+N6PBET+LnoFFBRcrK
hBgTi1VIuM/+Kwv3Mf6GLa3g9WI8vl9qhoE0Cymf8/8utXUvURK29HeFwhPKkeBd
DTlfHiZM6Fo/ymucFAMUdwN0Aalo5wzT9eshW1VttrDUe+v3bqPyymbmPSmZrLbt
WM1cdKqYskP2WOvm92s/HQZEdy0aohF+sGYlSvM75d6EMVEH7Y+5OgIslBcD/cgZ
5le9prjTSI6WEsV34CVdo9U8XNdFJjBZsUnNzqHixvev2fSFC9Ax/yu9XQZvmVxb
hz04pxmOVm+Mfxy78T29cIH1CMnNwOc2fH9uWi6iqD9k+79/EMeIg9fYUKLzXTCi
oBOfQNsdaQB4f63gy458ZhevA4wm14EgacrZEuCggLwh8KgwzpCROExzmFxc0e63
Om6M0hcD1B+G31GTr5PARHfINKi6osHatrYzgGoOYDkq2Jn0N/1Gy0a6+X/K1zRp
4/aiYODlD2vXiI4rLqbdQ+td1PVCB9Xrr4MXs+HGBn1YfNGhBgzNWjYDCEiVVgxY
FVj0Vc8CaaJD9I60oVG0KUKOGhDeqkAeKpdLqHWkAzILagpndh5hv1tH2LkmxVya
ojMdbD2Zd856Sb18PduFiBC3A0+uQDjuyZIZx/E3Ph1AX06bx3NeUzLKf38wq6eF
duBHivdpBO6osjG/WdpN26lmX58P2h12W1BzxmzbFaqWQjs+dzt7+9R6hER6b4i/
Apn/kqmPzUoJQEFR86z80d2hQO0AQpgS8jSYHEPZlne7h2lznyu7NuIRDTkf1yRi
v0cpDmCKkM8YoZgH5ioPffYmbvjrzVCxFv/fbPGsNeztc5PBZ/fFH3JvvysyfAB8
+zSONiDR/dZjOqKdJJURQOQ2yXUV/SU4WSuB+cyB5lnjrqFCKnyuJIeHLsXd3d8+
ud6iyVLDyA0inrmtxZVMCMqZyxpfmHom+ekECIxNr6v/MBC0TEdLhGAvYM0Q2SPV
0KedQt/bCbJIbup6PRIY/7z06WcDgJUACiSLiRstbWqoRBxznsI9Kw/ZudcZsBrz
8p+SD/qeFONzNDVSDsGV5vAmB6/ZDDQTMFLmapyaXD0cnik8F4h7PHK8MvZtBoBt
A7Sie9MYcdlGc3PQ74Ld2b15x8DW+dnMX3BjMzsqAbB+x2Qoka9nVpJF0fRwdzLY
hd4b1wzGoJzKiDGcSDGqvi/+/aiTXUY1i7yK3/uu7lXdoZrISFWYvYbMyiqsYmBF
dx42PtX2DCwpSotSgXMalAbFn5QW4CfPE3sGLlyVN9+1BZQdm1mFkQZOiDnceKc7
SBjch0FCZKMR1s/HE7FvPjYP5Qu78GRBQ//aqK4wBmfm52Kax7x6R+3Fc8VGIyEd
tU2vNaYxYpYVPd269A5DP6rrwHdGtPvtEs3lOEpNqNuI+/fl9JJqZPQNGXqlFILA
WtRMT995Jdf6OQz1ntMQqA2lB15205tIMYHEJJn2W8Q2/isch7SPbdepEuTKc7y9
hZ81ZEsQ4NiPCP7tCLRUQZoPUubJVPy5yjHXBlCx3VAOWRG2EulsYgt/McxvQyZm
zRu1UmRx3aMqzLI0ZDyP8pkQfQbE2Kq9EIEQ02AYQLWO2JZ4Z42y88U77YRg3GYC
EIpHT97+LHpTB8CVCb8tUDt4H0vEB8+vkJmN+jAOphnSnkKR+puEV1Oflxrn6LWi
1m/8IMzgr6DiQul9jOZL5B/3LXQWOENQLam+vwoCtXCGqvN2Ab8sP5bcyk8gEPFF
zvPyVoNEpJrHRpO9Fo5vIqf59xxPz+cbooboaWDCXfTLZ2ryuEMB3/fpc1e6Syv6
WtNUZafHe4KvaiXLb5kHSNbnPOOLU8xHGpZgDeTddeLBBqc+kUdEg4FzMeJhLdxE
MaAlLVeKQNONY0TRvkWzajZYGUs5waBcaDCRh6tkFqA9MDzTPjLBsce7mEO/UjVQ
RuV4n2Zdzqmu5ByYYV6DM+dVF5qbTxdF446ZXOpVBHiQ1y0cMb2jXK9bFIDArMB8
Rx1BhDvjlfpscM+jyUTDjkUh1HWkHahA6EcBCZBCkkz9LKDsktEeMIloI0AVruh/
3rYFXMeoZr8Hyy+B81xrdCsw65rSQhek2F2e2+TxqmtltqlVINuw5Uh889TkVeYx
25avVuYJIJstL8YN0yOghChqY7I2BTv14RppC20SX09EaO/eOzdL+BHvMXc+4Yzb
DA8MNSBRaLUHhozPMWy5ckgGEDP4uIEXA+tiyo5BIEqluoHiW0Ufv210seN90++N
3rgCaLt8OckgwTcISicyK3Ix8qIHsy8t4NgAAU0wzmKBFxBMiXV4J2HLoo3QyC1d
mwng37mbJI0N1at+4qaxqkcJyOJuIX3UWGg5NnQog7uSNcTYFRYTCVSuL3FjpQTQ
MSXrD5Lw/Qa2UhrIqi5aTohi1xoE3BonLIZbQZVxuYXyGay84/gdxLEPK+JM63eZ
R0E82KDTFbkz+OWzbBn694DuT6FXrWCsSfHz027RIJrwPTzVXntfpoWP/+299vgu
30sSiqmb3R3zHDBxFDMkUgRwSJ8vgTdEoNU7J1R4Qir3LApFERXcjnqEWUlia8ro
7upaxi5sZ6ns3+wWtA8MS3DJfRf30iHqqRw1UKuM8w3JeyJho5O8ByxsFhasAHRQ
Fk7OK3XRixUFFmEM6+2PWXSp/vZ9Zjkf1hLf6yj/CBpTGPYDZusp6SiKSxeibsth
+7ge8VlWReY5Et3YZGw1Y125VTj4J4jfXTBCdMH0kmQbRKXaFAZzhpKhwV28AFaw
pXW8xJS31QCpiMQK/koeb7eqQa0ryuQq+dZjTFlTWC2Uf+x2BZEG9E5GLucu9/Kn
gH1Bak+Yp7ZJ8KITAu4fbdM9awYWuFd86CyEwPkiNcxxhhR9yA0B1XoAMc/z+FZS
LKzr4dLj8fWESfX0A6rBHHtEs3291uZU80Qm8+UIoqrdIuq3jHQdd2VlgRDIcc6r
fsCBC66Ed6G02kEIH2URr7CrU+sKcz1F7QVyltwgQn7+eu42N9RyMwVK4FDRdMm9
XwqzNKrUTbrRRg17j/Dv6HVSXNd3317MLpk2dOKn/4D7Odah8ZhEhxReFtAw8RAg
FWgd3eP7+7OUu5MDxEGjVPwfkoX5DJNRdr3Tx33vsi9bmfaGo3VRbBJ9Jnh1DKy3
QNwjuOUn7XAtt97WlzPUe/4+7L45EyqvPOfrkjb9pNe2ZeaKHXEE6ItRsWyicLDN
wzZ3ZGmrdUWC8mMm5DWRJ6KeBXch3JrJgrwonrRKgmNbVsXae9FyG6D7aNC9pb2e
E0jCJuCKScsmu2ng29M6lka2HTXBzNXXD6ow7HnwGvY+2BlSOifG4KrpN98K0yzh
AyJE9qcUXs1zds2Wu0mtejYyrQfcDng8ixGelYWH9i0BPKzQRx/jghM3quKucQmS
HDmLcDiq29aBg/zcrJDyGz0GFWHjxMlPJGrqSqtWXmfbkQuwknoh59YQPUQzEkOP
+XqKlhaKUrJTF7fyKhck2WNNELjaUW782JUbQsHN8s4gYih2TAzoG9gKcJ1OgM0A
B33SU6mpvyN/RLY3UWT/GicT7YyF+uf469fCenYUu01dt4LFFssLAl6mrEatI+PD
Mc3h2RRKVnJs7SegPVSDune12b8OCbqVNO6Ln8TPM29Nvqu2Y3iomEz2WELs9NXg
14/L/otJmpkAbF9JEDYLBlv95Lv8r/MkLKF5+1vO5ZkfxjSXHNYJT7XsdH9vhhGO
J+lW/p/qI675pqT8Jj7isZ/4jW9Y0WzwwvBuJu72JfY2TH1R3gNtQ/IoAPNa0ivm
sY24o+0dKl04ExptSfH6GPsfOk4Qi2a4JlmSsELVGkyYdRo/znN8id8GR+dSXSUG
n5h+nHZaHfGUpS1x17qJLn13O+lwdbMfhVRMylGDZ5Hhipk2xSxJjkri01BdpImz
fJBfxI3nk10fPSBc6AFn2Z7SdNTIVtsi1Pp7s0AgNtW4tbUrdH7H2fDIbhpvnMsf
kftb/dVI3eUdzA7WrtVn81GkzyFfhyuDJikGgBpdrGpJw4HE7Mot7BjygAwd6xNF
6OuFO93boN8Ku9a91O06LwNylXPKditDGUAXtyQbsaTT/HAMUe40+5nz1/nr+x0g
B7mZ6ASYMZthkjCCeyd8FCpcH56i20jndSsoAt+usFdLm2NyBheRUjBMFJK2pxr9
any/9NzzccyEw6rNY3y+3ICyT1Z+cOFFQRFFCLswNgeza3vLHkZSROCc78783VGI
On+EyySlBFBR+6OeJ44VC6QkOv0y80i71fUtVHFzU+GNEqxsyWRjH23Sl8asyQwJ
R3OjT3TO2iBiK/7o1A3L6QQ+Ii6xlV3aO0ml4t2nwcyjd0g3+ii9870tzfJUgeA4
axUT6YCpo5jzbLjme9zyUeplX7sfFZs4GcH1E8T31BBavQ1Thj8xYIrarfMNKSw9
ZJUZdeUEVYc8dbZYFSomF26G+qO2cCcN7hbheSIBCjlAzffh3eXu/Xl2LFDMZSry
EIuYM0S7rhz1zJx+NegH3UnNe0d30h2YqWatpu0oDnqDv+TJDGJq3uQPgmhXrAeQ
J/ejpqDe3ruYwhUaFPkReNx02out0ZFMPv1CCgtPfYkbgiXi2s/YyBGAoIFkLBRO
tjRyNjzO7cwdInU54Ablg7geEYXfaCeDjZp0AVV0wl2eGGbuWXIo5RsofVuRHKoO
EDFbkGV8DD55vZ4IaoLk6lSTttttZfz19d1G7AiindZcqj5Gv1Tpvs9rdwJ2lcFr
JvsDjasMcgN5KV8+70F5GTg90rsNoFPiKPWzsUcNYCz3BS75APhfaoOh7FNcvLyS
PPUZY8GvE8uh6hhfbo1fxE8IqRufeKmlgqoepaZ2lgOsLPh+aw3L7Qs3WWLq1g8P
Q9MWK3geaQw8euCdQFA3efK/EQ6NBKsAOYtmh4tx167CXT0I2Zg9dBD6obwm7L0Q
Bo+FwXk9AYMW45Uw77mvEe6fIJcufRvXJEmlM5HW5BwCtE+s2czPpb84x0EWGItP
2dYdcQdYlwIM7wdUXQ15/V2KhzBijBW3OMaKLgHBEv54AG/XUr6IovyUZ8hrlNsy
Dyf12+T7E3OjTEwNBRvSneu4Z7Gf2WQIRajimu5eLNMC/InyJJvk1IDyrQNoxM/o
WLPrS3F1JN32Q+189whruFh7ivAthhluStwx/L4N9hjvwy3vx4ql63bkh2wmbnWj
vryUdaaPpnD8zodasj0LibJAJdZsRBhOY/xpR/pDWO3l+jrRYg1Bzgq3//U42VLh
vslG+pL01gb/5UFYY49pojdS95VdtrT5zlIbdmtMAPoMAKtimcudyt1YZgGUHpVf
LiOm0Ih8nwWHeRO+vT+2vvNLm2aYsLHqDIO0fKIAlcjhiumTJCqWsjHmoZNZOapf
DHE0Cei2EU10hcnsdsL21R5BjNXBmTqoBLgnfjykXxtowifpr+NPFEexPN3DRvFl
17Azsn1E7fcdR1uM6Cv4fkJBQHNVLKbAULiNO7xjzPwL0Xgve1dtW9iFi4ARWup8
4dwA98yGdEys/08CiPF3+pc9fyzEYwUfA/HSpQyMEpanyx2cxScjCxl8h+BfCeyG
joWo7zJcPbRD0tMs+E6WX13Eeg4Z9TyMoGOBMSw8o5RaLtp4E4j7ySoS0vlEixJh
9qMtmvT5MBrFp3RvlBfxyYS+EjXZwZYFOiB7aLrbSRXnyQfI1IR5IDy1WXlAM3vq
hKYnvtDiX61c0avyWWRSrPMeVRPN1gCwBKpL0p7wmoF2PZgC9NofT5TP7AcCQgWQ
h8rRYox9z8fmVOwFgEwhAHtN/2jFkV6CDErrR/PBlbZXAFCnpL+mNpaytxz7LeWi
FChQIHE3sTJa0VAm3Nc/Blb4ObDW0A5wr5xm5xfLyRmxqwBf4Gix4UZaeDh4/SJT
3rzhl6J3sS0EbxY5TPUkFFq3gi/r3tEr/Wb78J04pjT0Ugs10Z9zVPnQbrWCulVm
xKyqKJ97rd/7b6Yus/Nr/9t2ESiuQl1zro3EjOrmQW7lh1PemYcaFKOFPaJeMzkH
cJ9HZRfxzOdtYWnkwcDzIGVBen/7qwQFSbvpnkXqqUX21XzBQGWuNfxTcq/hr9UA
J+N/HrFJkaY+ZYbJLlXz7pV9dXmJ6LIaJ/acm0U+SnVZ8yD05IHf/2yaAtzhlVDc
2kLzGCJ3Jd5pXMz2aO4PO/8NOhnwCOmQFX4qOSAHobLjYRJ1HQbV5zaPwz+/fdxB
BTnDj9aPHs/5hbGEOk3W28mebuKYzo3+T7Wt9rCs/5iGatNX2Gy83nfkMVoFtm+p
YtzYO70is8lGVeGoTvzJI7ldnJfo11R8B2ncWrk8c8WKllGh3YCU3MbJQb5Zanea
V6VlacywHXR5gMgAVMAkcDpgT7lvvJO/WGP392sEROqgrMrSNm1NQuple7rM2DYX
qy1cc2YnSt5IsRfFKeTZ4hSkHs5+JUMeBn7WkM26y6ZB8Y9kGJmhOX2QBIx9q7OX
RzT0jRCvlHNmeAa65gq9mHBTyhZThznjmYaOCVN4rk5cOeUOkW6EDu/sBdraUiQm
t+HtDJA6dpAS1zN0j4KbecrXmwsQbmQl4Uj+cyTSrOY2w76fFKd+gizRwtF+5GLK
JoD90AbZ9MHj72PUCzPecdsdvumnHPAr4//zOEnpQHDvYvTDrfeQMLf7NXq6o0sX
armBRgOP47t3LwZWnlfRV6pxgjSycg1BTbjhJnAe220z3kqrO1QGmkQprdGLROB/
VVQPUq+47TQlsQDCmsarBUPKz/AzxwlLeucwLzKeqqPFhi7EzVD/mpTUsSiXDIVH
fbGmpZK48rsbOFZgZkB7xWY0n9Nnp4gRT30AHsIFE5u6ewjkYBlA2LrVN0NJIeOn
i8pWzeEcI/J3w8fhkf9DKQgIqf4+qOezJFuo0lWFL5lMkX907rHK8Uqb0zE11+sT
lhHDsYcddQMxXqj0rtb17nsShkN5vHGPEcXRvoj8QSZS8bESFHHff94qWK8bxGvh
XXrvw/znVQa9ArReUlxpiKXgoR7EkohTEGeuAy95lT6oaHyQGhgvppyskqkJW4dI
hVqa0iphKLsY64Bfr9a5kH4Nh1SherChoItquCK7mFQXKcYXWJJudYwSFdwnq/lN
1sbHzlxfe4SYZs70k9fTvRdL/Exzv/lrpFhFv6P3xc6ukNzv/dV4Mjwd4pqNCdVQ
`pragma protect end_protected
